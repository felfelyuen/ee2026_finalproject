// Revision:`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 11.04.2025 00:50:31
// Design Name: 
// Module Name: start_screen
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 

// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module felix_start_screen(
    input [6:0] x,
    input [5:0] y,
    output reg [15:0] start_screen_data
    );
    
    always @ (*) begin
        if ((y == 6 && ((x >= 40 && x <= 44) || (x >= 49 && x <= 52) || (x == 56 || x== 57 || x == 63 || x == 64) || (x >= 67 && x <= 71))) // "BOMB"
            || ((y >= 7 && y <= 15) && ((x == 40) || (x == 48) || (x == 53) || (x == 56) || (x == 64) || (x == 67)))
            || ((x >= 41 && x <= 44) && (y == 11 || y == 16))
            || (x == 45 && ((y >= 7 && y <= 10) || (y >= 12 && y <= 15)))
            || (y == 16 && (x == 40 || (x >= 49 && x <= 52) || (x >= 55 && x <= 57) || (x >= 63 && x <= 65) || (x >= 67 && x <= 71)))
            || (y == 7 && (x == 57 || x == 58 || x == 62 || x == 63 || x == 72))
            || (y == 8 && ((x >= 57 && x <= 59) || (x >= 61 && x <= 63) || x == 72))
            || (y == 9 && ((x >= 58 && x <= 62) || x == 72))
            || (y == 10 && ((x >= 59 && x <= 61) || x == 72))
            || (y == 11 && ((x == 60) || (x >= 68 && x <= 71)))
            || (x == 72 && ((y >= 12 && y <= 15)))
            || (x == 46 && y >= 21 && y <= 27) //"GO"
            || (x == 47 && ((y >= 20 && y <= 21) || (y >= 27 && y <= 28)))
            || ((y == 19 || y == 29) && ((x >= 48 && x <= 52) || (x >= 57 && x <= 60)))
            || (x == 52 && (y == 20 || (y >= 24 && y <= 28)))
            || ((y >= 20 && y <= 28) && (x == 56 || x == 61))
            || (y == 24 && (x == 51 || x == 53))
            || ((y >= 33 && y <= 41) && (x == 40 || x == 48 || x == 53 || x == 56 || x == 61 || x == 64 || x == 72)) //"BOOM!"
            || ((x >= 41 && x <= 44) && (y == 32 || y == 37 || y == 42))
            || (x == 45 && ((y >= 33 && y <= 36) || (y >= 38 && y <= 41)))
            || (x == 40 && (y == 32 || y == 42))
            || (y == 32 && ((x >= 49 && x <= 52) || (x >= 57 && x <= 60) || (x >= 64 && x <= 65) || (x >= 71 && x <= 72)))
            || (y == 42 && ((x >= 49 && x <= 52) || (x >= 57 && x <= 60) || (x >= 63 && x <= 65) || (x >= 71 && x <= 73) || (x == 76)))
            || ((y >= 32 && y <= 34) && (x == 65 || x == 71))
            || ((y >= 33 && y <= 35) && (x == 66 || x == 70))
            || ((y >= 34 && y <= 36) && (x == 67 || x == 69))
            || ((y >= 34 && y <= 36) && (x == 68))
            || (x == 76 && y >= 32 && y <= 39)) begin
            start_screen_data = 16'b11111_111111_11111;
        end else if (x == 3 || x == 4) begin
            start_screen_data = 16'b11111_100000_01101; //pink wire
        end else if (x == 9 || x == 10) begin
            start_screen_data = 16'b11111_000000_00000; //red wire
        end else if (x == 15 || x == 16) begin
            start_screen_data = 16'b00000_000000_11111; //blue wire
        end else if (x == 21 || x == 22) begin
            start_screen_data = 16'b11111_101001_00000; //orange wire
        end else if (x == 27 || x == 28) begin
            start_screen_data = 16'b00000_111111_00000; //green wire
        end else begin
            start_screen_data = 16'b00000_000000_00000; //black background
        end
    end
    
endmodule