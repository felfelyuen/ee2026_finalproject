// Revision:`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 11.04.2025 00:50:31
// Design Name: 
// Module Name: start_screen
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 

// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module felix_start_screen(
    input [6:0] x, //column number
    input [5:0] y, //row number
    output reg [15:0] olede
    );
    
    always @ (*) begin
        olede = 16'h0000;
        //black background
        if (x >= 6 & x <= 86 & y >= 12 & y <= 53) begin
            olede = 16'hFFC2; //yellow sign
        end
        
        if (((x == 27 | x == 28) & (y <= 63 & y >= 58)) |
         ((x >= 27 & x <= 95 & y >= 58 & y <= 59 ))) begin
            olede = 16'hFC0D; //pink wire
        end 
        else if ( (x >= 21 & x <= 22 & y <= 63 & y >= 54) | 
        (x >= 21 & x <= 95 & y >= 54 & y <= 55) |
        (x >= 90 & x <= 95 & y >= 18 & y <= 19) | 
        (x >= 87 & x <= 89 & y >= 17 & y <= 18) | 
        (x >= 74 & x <= 76 & y >= 9 & y <= 11) |
        (x >= 73 & x <= 75 & y >= 7 & y <= 8) |
        (x >= 73 & x <= 74 & y >= 5 & y <= 6) |
        (x >= 72 & x <= 73 & y <= 5)) begin
            olede = 16'hF800; // red wire
        end 
        else if ((x >= 15 & x <= 16 & y <= 63 & y >= 50) | 
        (x >= 15 & x <= 95 & y <= 51 & y >= 50) | 
        (x >= 84 & x <= 95 & y <= 25 & y >= 24) | 
        (x >= 83 & x <= 84 & y <= 24 & y >= 22) | 
        (x >= 82 & x <= 83 & y <= 23 & y >= 20) |
        (x >= 81 & x <= 82 & y <= 21 & y >= 15) |
        (x >= 82 & x <= 83 & y <= 14)) begin
            olede = 16'h001F; // blue wire
        end
        else if ((x >= 9 & x <= 10 & y <= 63 & y >= 46) | 
        (x >= 9 & x <= 95 & y <= 47 & y >= 46) |
        (x == 22 & y == 39) |  
        (x >= 21 & x <= 23 & y == 38) |
        (x >= 20 & x <= 24 & y == 37) |
        (x >= 19 & x <= 25 & y == 36) |
        (x >= 18 & x <= 26 & y == 35) |
        (x >= 17 & x <= 27 & y == 34) |
        (x >= 16 & x <= 28 & y == 33) |
        (x >= 15 & x <= 29 & y == 32) |
        (x >= 14 & x <= 30 & y == 31) |
        (x >= 13 & x <= 31 & y == 30) |
        (x >= 12 & x <= 32 & y == 29) |
        (x >= 13 & x <= 31 & y == 28) |
        (x >= 14 & x <= 30 & y == 27) |
        (x >= 15 & x <= 29 & y == 26) |
        (x >= 16 & x <= 28 & y == 25) |
        (x >= 17 & x <= 27 & y == 24) |
        (x >= 18 & x <= 26 & y == 23) |
        (x >= 19 & x <= 25 & y == 22) |
        (x >= 20 & x <= 24 & y == 21) |
        (x >= 21 & x <= 23 & y == 20) |
        (x == 22 & y == 19)) begin
            olede = 16'hFD20; //orange bits
        end
        else if ((x >= 3 & x <= 4 & y <= 63 & y >= 42) | 
        (x >= 3 & x <= 95 & y <= 43 & y >= 42) |
        (x >= 4 & x <= 7 & y <= 24 & y >= 23) |
        (x >= 7 & x <= 9 & y <= 23 & y >= 22) |
        (x >= 9 & x <= 11 & y <= 22 & y >= 21) |
        (x >= 10 & x <= 12 & y <= 20) |
        (x >= 11 & x <= 12 & y <= 20 & y >= 18) |
        (x >= 12 & x <= 13 & y <= 18 & y >= 15)) begin
            olede = 16'h07E0; //green bits
        end
        else if ((x == 22 & y == 40) |
        ((x == 21 | x == 23) & y == 39) |  
        ((x == 20 | x == 24) & y == 38) |
        ((x == 19 | x == 25) & y == 37) |
        ((x == 18 | x == 26) & y == 36) |
        ((x == 17 | x == 27 |( x >= 70 & x <= 74)| (x >= 61 & x <= 68) | (x >= 56 & x <= 59) | (x >= 46 & x <= 54) | x == 41 | x == 43 | x == 44) & y == 35) |
        ((x == 16 | x == 28) & y == 34) |
        ((x == 15 | x == 29) & y == 33) |
        ((x == 14 | x == 30) & y == 32) |
        ((x == 13 | x == 31) & y == 31) |
        ((x == 12 | x == 32) & y == 30) |
        ((x == 11 | x == 33 | x == 55 | x == 48 | x == 42) & y == 29) |
        ((x == 12 | x == 32 | x == 54 | x == 47) & y == 28) |
        ((x == 13 | x == 31) & y == 27) |
        ((x == 14 | x == 30) & y == 26) |
        ((x == 15 | x == 29) & y == 25) |
        ((x == 16 | x == 28) & y == 24) |
        ((x == 17 | x == 27 | (x >= 62 & x <= 74) | (x >= 52 & x <= 60) | (x >= 48 & x <= 50) | x == 46 | (x >= 41 & x <= 44)) & y == 23) |
        ((x == 18 | x == 26) & y == 22) |
        ((x == 19 | x == 25) & y == 21) |
        ((x == 20 | x == 24) & y == 20) |
        ((x == 21 | x == 23) & y == 19) |
        ((x == 20 | x == 22) & y == 20) |
        (x == 21 & y == 20) |
        (x == 74 & y <= 32 & y >= 28) |
        (x == 70 & y <= 32 & y >= 28) |
        (x == 72 & y <= 29 & y >= 27) |
        (x == 68 & y <= 31 & y >= 27) |
        (x == 64 & y <= 31 & y >= 27) |
        (x == 62 & y <= 31 & y >= 27) |
        (x == 58 & y <= 31 & y >= 30) |
        (x == 58 & y <= 28 & y >= 27) |
        (x == 56 & y <= 32 & y >= 27) |
        (x == 53 & y <= 32 & y >= 27) |
        (x == 51 & y <= 32 & y >= 27) |
        (x == 49 & y <= 32 & y >= 27) |
        (x == 46 & y <= 32 & y >= 27) |
        (x == 44 & y <= 31 & y >= 28) |
        (x == 41 & y <= 29 & y >= 28) |
        (x >= 65 & x <= 67 & y == 32) |
        (x >= 65 & x <= 67 & y == 28) |
        (x >= 59 & x <= 61 & y == 32) |
        (x >= 59 & x <= 61 & y == 28) |
        (x >= 41 & x <= 43 & y == 32) |
        (x >= 42 & x <= 43 & y == 27) |
        (x >= 59 & x <= 61 & y == 28) |
        (x >= 71 & x <= 73 & y == 27)) begin
        olede = 16'h0000; //black bits
        end
        
        if ((x >= 21 & x <= 23 & y <= 35 & y >= 28) |
        (x >= 21 & x <= 23 & y <= 25 & y >= 23)) begin
        olede = 16'h0000;
        end
        
    end
    
endmodule
