`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 04/12/2025 02:52:04 PM
// Design Name: 
// Module Name: picture_converter
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module picture_converter(
input CLK,
input [12:0] pixel_index, 
output reg [15:0] oled_data
    );
    
    always @(posedge CLK) begin
    if (pixel_index == 0) oled_data = 16'b0011101010000100;
    else if (pixel_index == 1 || pixel_index == 99 || pixel_index == 102 || pixel_index == 613 || pixel_index == 924 || pixel_index == 1582) oled_data = 16'b0100001011000101;
    else if (pixel_index == 2 || pixel_index == 3841) oled_data = 16'b0011101010000101;
    else if (pixel_index == 3 || pixel_index == 104 || pixel_index == 2579) oled_data = 16'b0100001100000100;
    else if (pixel_index == 4 || pixel_index == 395 || pixel_index == 1842) oled_data = 16'b0101001100000110;
    else if (pixel_index == 5 || pixel_index == 105 || pixel_index == 296) oled_data = 16'b0100101100000110;
    else if (((pixel_index >= 6) && (pixel_index <= 7)) || pixel_index == 926 || pixel_index == 1004 || pixel_index == 1207) oled_data = 16'b0100001010000101;
    else if (pixel_index == 8 || pixel_index == 616 || pixel_index == 1001 || pixel_index == 1684 || pixel_index == 2843) oled_data = 16'b0100101011000101;
    else if (pixel_index == 9) oled_data = 16'b0100101011001000;
    else if (pixel_index == 10 || pixel_index == 1306 || pixel_index == 2734 || pixel_index == 3556) oled_data = 16'b0101001100001001;
    else if (pixel_index == 11 || pixel_index == 2072) oled_data = 16'b0101001100001010;
    else if (pixel_index == 12) oled_data = 16'b0100101011001010;
    else if (pixel_index == 13 || pixel_index == 252 || pixel_index == 592 || pixel_index == 5251) oled_data = 16'b0100001011001100;
    else if (pixel_index == 14) oled_data = 16'b0011101010001101;
    else if (pixel_index == 15 || ((pixel_index >= 227) && (pixel_index <= 228)) || pixel_index == 253) oled_data = 16'b0011001011001110;
    else if (pixel_index == 16 || pixel_index == 2496) oled_data = 16'b0011001010001111;
    else if (pixel_index == 17) oled_data = 16'b0010101001010001;
    else if (pixel_index == 18 || pixel_index == 21 || pixel_index == 32 || pixel_index == 116) oled_data = 16'b0010001000010001;
    else if (pixel_index == 19 || pixel_index == 48 || pixel_index == 52 || pixel_index == 63 || pixel_index == 115 || pixel_index == 127 || pixel_index == 132 || pixel_index == 258) oled_data = 16'b0001101000010001;
    else if (pixel_index == 20) oled_data = 16'b0010001000010010;
    else if (pixel_index == 22 || pixel_index == 119 || pixel_index == 257) oled_data = 16'b0001101000010010;
    else if (pixel_index == 23 || pixel_index == 126 || pixel_index == 162 || pixel_index == 356 || pixel_index == 364 || pixel_index == 372 || pixel_index == 375 || pixel_index == 466 || pixel_index == 471) oled_data = 16'b0001001000010010;
    else if (pixel_index == 24 || pixel_index == 36 || pixel_index == 43 || pixel_index == 138 || pixel_index == 171 || pixel_index == 260 || pixel_index == 275 || pixel_index == 278) oled_data = 16'b0000100111010010;
    else if (pixel_index == 25 || pixel_index == 68 || pixel_index == 122 || pixel_index == 140 || ((pixel_index >= 164) && (pixel_index <= 165)) || pixel_index == 167 || pixel_index == 237 || pixel_index == 261 || pixel_index == 279) oled_data = 16'b0000000111010010;
    else if (((pixel_index >= 26) && (pixel_index <= 28)) || pixel_index == 39 || pixel_index == 44 || pixel_index == 46 || pixel_index == 137 || pixel_index == 150 || pixel_index == 166) oled_data = 16'b0000000110010010;
    else if (pixel_index == 29 || pixel_index == 31 || pixel_index == 61 || pixel_index == 134 || pixel_index == 161) oled_data = 16'b0001000111010001;
    else if (pixel_index == 30) oled_data = 16'b0001000110010001;
    else if (pixel_index == 33) oled_data = 16'b0001100111010001;
    else if (pixel_index == 34 || pixel_index == 76 || pixel_index == 81 || pixel_index == 86 || pixel_index == 88 || pixel_index == 90 || pixel_index == 93 || ((pixel_index >= 169) && (pixel_index <= 170)) || pixel_index == 176 || pixel_index == 186 || pixel_index == 188 || pixel_index == 280) oled_data = 16'b0000100111010000;
    else if (pixel_index == 35 || pixel_index == 53 || pixel_index == 163 || ((pixel_index >= 264) && (pixel_index <= 265)) || pixel_index == 272 || ((pixel_index >= 282) && (pixel_index <= 285)) || pixel_index == 370 || pixel_index == 564) oled_data = 16'b0000101000010001;
    else if (((pixel_index >= 37) && (pixel_index <= 38)) || pixel_index == 56 || pixel_index == 65 || pixel_index == 67 || pixel_index == 69 || pixel_index == 72 || pixel_index == 87 || pixel_index == 89 || pixel_index == 135 || pixel_index == 143 || pixel_index == 152 || pixel_index == 172 || ((pixel_index >= 179) && (pixel_index <= 184)) || ((pixel_index >= 270) && (pixel_index <= 271)) || pixel_index == 274) oled_data = 16'b0000100111010001;
    else if (pixel_index == 40) oled_data = 16'b0000100110010001;
    else if (((pixel_index >= 41) && (pixel_index <= 42)) || pixel_index == 54 || ((pixel_index >= 70) && (pixel_index <= 71)) || pixel_index == 151) oled_data = 16'b0000000110010001;
    else if (pixel_index == 45 || pixel_index == 66) oled_data = 16'b0000000111010001;
    else if (pixel_index == 47 || pixel_index == 58 || pixel_index == 185 || (pixel_index >= 189) && (pixel_index <= 190)) oled_data = 16'b0001000111010000;
    else if (pixel_index == 49) oled_data = 16'b0100101100010100;
    else if (pixel_index == 50 || pixel_index == 221 || pixel_index == 432 || pixel_index == 583) oled_data = 16'b0011001011010010;
    else if (pixel_index == 51) oled_data = 16'b0010001000010011;
    else if (pixel_index == 55 || pixel_index == 74 || pixel_index == 79) oled_data = 16'b0000000110010000;
    else if (pixel_index == 57 || pixel_index == 142) oled_data = 16'b0000000110010011;
    else if (pixel_index == 59 || pixel_index == 117 || (pixel_index >= 211) && (pixel_index <= 212)) oled_data = 16'b0010001001010001;
    else if (pixel_index == 60 || pixel_index == 131 || pixel_index == 160 || (pixel_index >= 498) && (pixel_index <= 499)) oled_data = 16'b0010001001010000;
    else if (pixel_index == 62) oled_data = 16'b0001001000001111;
    else if (pixel_index == 64 || pixel_index == 191) oled_data = 16'b0001001000010000;
    else if (pixel_index == 73 || pixel_index == 77) oled_data = 16'b0000100110001111;
    else if (pixel_index == 75 || pixel_index == 82 || pixel_index == 85) oled_data = 16'b0000100110010000;
    else if (pixel_index == 78 || pixel_index == 91) oled_data = 16'b0000000110001111;
    else if (pixel_index == 80 || pixel_index == 92 || pixel_index == 168 || ((pixel_index >= 173) && (pixel_index <= 175)) || ((pixel_index >= 177) && (pixel_index <= 178)) || pixel_index == 187) oled_data = 16'b0000000111010000;
    else if (pixel_index == 83 || pixel_index == 94) oled_data = 16'b0001000111001111;
    else if (pixel_index == 84 || pixel_index == 95) oled_data = 16'b0000100111001111;
    else if (pixel_index == 96 || pixel_index == 519 || pixel_index == 1095) oled_data = 16'b0011001011000110;
    else if (((pixel_index >= 97) && (pixel_index <= 98)) || ((pixel_index >= 198) && (pixel_index <= 199)) || pixel_index == 640) oled_data = 16'b0100001011000110;
    else if (((pixel_index >= 100) && (pixel_index <= 101)) || pixel_index == 1494) oled_data = 16'b0100101011000110;
    else if (pixel_index == 103 || pixel_index == 711) oled_data = 16'b0100001011000100;
    else if (pixel_index == 106 || pixel_index == 540 || pixel_index == 908 || pixel_index == 3555) oled_data = 16'b0100101100000111;
    else if (pixel_index == 107 || pixel_index == 392) oled_data = 16'b0100101011001001;
    else if (pixel_index == 108) oled_data = 16'b0100001011001010;
    else if (pixel_index == 109 || pixel_index == 4080) oled_data = 16'b0011101011001100;
    else if (pixel_index == 110 || pixel_index == 2882) oled_data = 16'b0011001010001101;
    else if (pixel_index == 111 || pixel_index == 207 || pixel_index == 254 || pixel_index == 303 || pixel_index == 521) oled_data = 16'b0010101010001101;
    else if (pixel_index == 112 || pixel_index == 225) oled_data = 16'b0010001010001110;
    else if (pixel_index == 113 || (pixel_index >= 208) && (pixel_index <= 209)) oled_data = 16'b0010001001001111;
    else if (pixel_index == 114) oled_data = 16'b0010001000010000;
    else if (pixel_index == 118) oled_data = 16'b0010001001010010;
    else if (pixel_index == 120 || pixel_index == 139 || pixel_index == 232 || ((pixel_index >= 235) && (pixel_index <= 236)) || pixel_index == 239 || ((pixel_index >= 246) && (pixel_index <= 247)) || pixel_index == 263 || pixel_index == 266 || pixel_index == 268 || pixel_index == 333 || pixel_index == 361 || pixel_index == 363 || pixel_index == 365 || pixel_index == 374 || ((pixel_index >= 376) && (pixel_index <= 378)) || ((pixel_index >= 380) && (pixel_index <= 382)) || pixel_index == 430 || ((pixel_index >= 467) && (pixel_index <= 468)) || pixel_index == 472) oled_data = 16'b0000101000010010;
    else if (pixel_index == 121 || pixel_index == 262 || pixel_index == 379 || pixel_index == 457 || pixel_index == 459 || pixel_index == 551) oled_data = 16'b0000001000010010;
    else if (pixel_index == 123 || pixel_index == 141 || pixel_index == 217 || pixel_index == 234 || pixel_index == 267) oled_data = 16'b0000000111010011;
    else if ((pixel_index >= 124) && (pixel_index <= 125)) oled_data = 16'b0001000111010010;
    else if (pixel_index == 128 || pixel_index == 210 || pixel_index == 355) oled_data = 16'b0001101001010001;
    else if (pixel_index == 129) oled_data = 16'b0001101000010000;
    else if (pixel_index == 130 || pixel_index == 230 || pixel_index == 305 || pixel_index == 401) oled_data = 16'b0001101001001110;
    else if (pixel_index == 133 || pixel_index == 286) oled_data = 16'b0001001000010001;
    else if (pixel_index == 136 || pixel_index == 153) oled_data = 16'b0000100110010010;
    else if (pixel_index == 144) oled_data = 16'b0011101100010001;
    else if (pixel_index == 145 || pixel_index == 1926 || pixel_index == 3134) oled_data = 16'b0111010010110010;
    else if (pixel_index == 146) oled_data = 16'b0101001110010000;
    else if (pixel_index == 147) oled_data = 16'b0100001011010010;
    else if (pixel_index == 148 || pixel_index == 689) oled_data = 16'b0011001100010001;
    else if (pixel_index == 149 || pixel_index == 451 || pixel_index == 837) oled_data = 16'b0001101010010010;
    else if (pixel_index == 154 || pixel_index == 304 || pixel_index == 400) oled_data = 16'b0010101010001110;
    else if (pixel_index == 155 || pixel_index == 2264 || pixel_index == 5171 || pixel_index == 5176) oled_data = 16'b0100101100010000;
    else if (pixel_index == 156) oled_data = 16'b0011101011001111;
    else if (pixel_index == 157 || pixel_index == 226) oled_data = 16'b0010101010001111;
    else if (pixel_index == 158) oled_data = 16'b0010101001010000;
    else if (pixel_index == 159) oled_data = 16'b0011001001010001;
    else if (pixel_index == 192) oled_data = 16'b0010101010001010;
    else if (pixel_index == 193 || pixel_index == 289) oled_data = 16'b0011101010001010;
    else if (pixel_index == 194 || pixel_index == 293) oled_data = 16'b0011001010001001;
    else if (pixel_index == 195) oled_data = 16'b0011001001001001;
    else if (pixel_index == 196 || pixel_index == 423) oled_data = 16'b0011001010000111;
    else if (pixel_index == 197) oled_data = 16'b0100001010000110;
    else if (pixel_index == 200 || pixel_index == 203 || pixel_index == 2478) oled_data = 16'b0101001100000101;
    else if (((pixel_index >= 201) && (pixel_index <= 202)) || pixel_index == 1409 || pixel_index == 1982 || pixel_index == 2574) oled_data = 16'b0101101101000101;
    else if (pixel_index == 204 || pixel_index == 1005 || pixel_index == 1017) oled_data = 16'b0101001100000111;
    else if (pixel_index == 205 || ((pixel_index >= 480) && (pixel_index <= 481)) || pixel_index == 811) oled_data = 16'b0100001100001001;
    else if (pixel_index == 206 || pixel_index == 386 || pixel_index == 3072 || pixel_index == 4272) oled_data = 16'b0011001011001100;
    else if (pixel_index == 213) oled_data = 16'b0010101001010010;
    else if (pixel_index == 214 || pixel_index == 310) oled_data = 16'b0010001010010010;
    else if (pixel_index == 215 || pixel_index == 367 || pixel_index == 475 || ((pixel_index >= 478) && (pixel_index <= 479)) || pixel_index == 571 || pixel_index == 575) oled_data = 16'b0001001001010010;
    else if (pixel_index == 216 || pixel_index == 312 || pixel_index == 331 || pixel_index == 335 || pixel_index == 653) oled_data = 16'b0000001000010011;
    else if (pixel_index == 218 || pixel_index == 314 || pixel_index == 334 || ((pixel_index >= 357) && (pixel_index <= 358)) || pixel_index == 371 || pixel_index == 373 || pixel_index == 431 || pixel_index == 462 || pixel_index == 473) oled_data = 16'b0000101000010011;
    else if (pixel_index == 219) oled_data = 16'b0001001000010011;
    else if (pixel_index == 220) oled_data = 16'b0010001001010011;
    else if (pixel_index == 222 || pixel_index == 388) oled_data = 16'b0010101010010000;
    else if (pixel_index == 223 || pixel_index == 387 || pixel_index == 485) oled_data = 16'b0010101011010000;
    else if (pixel_index == 224 || pixel_index == 352 || pixel_index == 486) oled_data = 16'b0011001011001111;
    else if (pixel_index == 229 || pixel_index == 291 || pixel_index == 826) oled_data = 16'b0010001010001101;
    else if (pixel_index == 231 || pixel_index == 306 || pixel_index == 402) oled_data = 16'b0001001001010000;
    else if (pixel_index == 233 || pixel_index == 238 || pixel_index == 313) oled_data = 16'b0000000111010100;
    else if (pixel_index == 240 || pixel_index == 585 || pixel_index == 1190 || pixel_index == 3073) oled_data = 16'b0100001101010000;
    else if (pixel_index == 241 || pixel_index == 1202) oled_data = 16'b1010111001101111;
    else if (pixel_index == 242 || pixel_index == 2241 || pixel_index == 2364) oled_data = 16'b0111110101101111;
    else if (pixel_index == 243) oled_data = 16'b0110110001010010;
    else if (pixel_index == 244) oled_data = 16'b0101101111010001;
    else if (pixel_index == 245 || pixel_index == 342) oled_data = 16'b0010101100010010;
    else if (pixel_index == 248 || pixel_index == 582 || pixel_index == 606) oled_data = 16'b0010101011010010;
    else if (pixel_index == 249) oled_data = 16'b0010101000010010;
    else if (pixel_index == 250) oled_data = 16'b0100101101001100;
    else if (pixel_index == 251 || pixel_index == 3459) oled_data = 16'b0101101110001010;
    else if (pixel_index == 255) oled_data = 16'b0011101011010000;
    else if (pixel_index == 256 || pixel_index == 328) oled_data = 16'b0010001010010000;
    else if (pixel_index == 259 || pixel_index == 281) oled_data = 16'b0000101000010000;
    else if (pixel_index == 269) oled_data = 16'b0000001000010001;
    else if (pixel_index == 273) oled_data = 16'b0000001000001111;
    else if (pixel_index == 276) oled_data = 16'b0000100110010011;
    else if (pixel_index == 277) oled_data = 16'b0000100111010011;
    else if (pixel_index == 287) oled_data = 16'b0001001001010001;
    else if (pixel_index == 288 || pixel_index == 398) oled_data = 16'b0100001011001001;
    else if (pixel_index == 290 || (pixel_index >= 1115) && (pixel_index <= 1116)) oled_data = 16'b0010101010001011;
    else if (pixel_index == 292 || pixel_index == 2881) oled_data = 16'b0011001011001011;
    else if (pixel_index == 294) oled_data = 16'b0011101001001000;
    else if (pixel_index == 295) oled_data = 16'b0011101010001000;
    else if (pixel_index == 297) oled_data = 16'b0100101110000100;
    else if (pixel_index == 298 || pixel_index == 2183 || pixel_index == 2475) oled_data = 16'b0101001101000011;
    else if (pixel_index == 299) oled_data = 16'b0100101100000100;
    else if (pixel_index == 300 || pixel_index == 1840) oled_data = 16'b0101001100000100;
    else if (pixel_index == 301) oled_data = 16'b0101001011000110;
    else if (pixel_index == 302 || pixel_index == 326 || pixel_index == 385) oled_data = 16'b0011101011001001;
    else if (pixel_index == 307 || pixel_index == 403) oled_data = 16'b0001001010010001;
    else if (pixel_index == 308) oled_data = 16'b0001101001010010;
    else if (pixel_index == 309) oled_data = 16'b0010001001010100;
    else if (pixel_index == 311 || pixel_index == 366 || pixel_index == 368 || pixel_index == 407 || pixel_index == 452 || pixel_index == 454 || pixel_index == 458 || pixel_index == 461 || pixel_index == 465 || ((pixel_index >= 469) && (pixel_index <= 470)) || pixel_index == 476 || pixel_index == 550 || pixel_index == 552 || pixel_index == 563 || pixel_index == 566 || pixel_index == 645) oled_data = 16'b0000101001010010;
    else if (pixel_index == 315 || pixel_index == 410) oled_data = 16'b0001101010010011;
    else if (pixel_index == 316 || pixel_index == 685 || pixel_index == 833) oled_data = 16'b0011001100010010;
    else if (pixel_index == 317 || pixel_index == 343 || pixel_index == 580) oled_data = 16'b0100101110010000;
    else if (pixel_index == 318) oled_data = 16'b0100001110001110;
    else if (pixel_index == 319 || pixel_index == 638) oled_data = 16'b0101001110001100;
    else if (pixel_index == 320 || pixel_index == 803 || pixel_index == 1891 || pixel_index == 2384) oled_data = 16'b0101001111001010;
    else if (pixel_index == 321) oled_data = 16'b0100101110001100;
    else if (pixel_index == 322) oled_data = 16'b0011101110001010;
    else if (pixel_index == 323 || pixel_index == 2386) oled_data = 16'b0011101110001001;
    else if (pixel_index == 324 || pixel_index == 2581) oled_data = 16'b0100001110001000;
    else if (pixel_index == 325 || pixel_index == 806 || pixel_index == 1421 || pixel_index == 2570) oled_data = 16'b0100101110000111;
    else if (pixel_index == 327 || pixel_index == 424 || pixel_index == 2497) oled_data = 16'b0011001010001100;
    else if (pixel_index == 329) oled_data = 16'b0000101000010100;
    else if (pixel_index == 330) oled_data = 16'b0000001000010101;
    else if (pixel_index == 332) oled_data = 16'b0000101010010001;
    else if (pixel_index == 336 || pixel_index == 581) oled_data = 16'b0011101101010010;
    else if (pixel_index == 337) oled_data = 16'b1100111011101100;
    else if (pixel_index == 338) oled_data = 16'b1000010111101011;
    else if (pixel_index == 339) oled_data = 16'b0110110100101101;
    else if (pixel_index == 340 || pixel_index == 2121) oled_data = 16'b0110010011101111;
    else if (pixel_index == 341 || pixel_index == 527) oled_data = 16'b0011101101010011;
    else if (pixel_index == 344 || pixel_index == 940 || pixel_index == 2063) oled_data = 16'b0111110011101111;
    else if (pixel_index == 345 || pixel_index == 3173) oled_data = 16'b0110101110001100;
    else if (pixel_index == 346 || pixel_index == 909 || pixel_index == 1653 || pixel_index == 2668 || pixel_index == 2821) oled_data = 16'b0110010000001001;
    else if (pixel_index == 347 || pixel_index == 1278 || pixel_index == 1577 || pixel_index == 1654 || pixel_index == 2383 || pixel_index == 2466 || pixel_index == 3324) oled_data = 16'b0110001111001001;
    else if (pixel_index == 348 || pixel_index == 489) oled_data = 16'b0100101100001010;
    else if (pixel_index == 349 || pixel_index == 482 || pixel_index == 589) oled_data = 16'b0100001100001100;
    else if (pixel_index == 350) oled_data = 16'b0011001100001011;
    else if (pixel_index == 351 || pixel_index == 496) oled_data = 16'b0011101011001101;
    else if (pixel_index == 353 || pixel_index == 450) oled_data = 16'b0011001010010001;
    else if (pixel_index == 354) oled_data = 16'b0010001010010001;
    else if (((pixel_index >= 359) && (pixel_index <= 360)) || pixel_index == 455) oled_data = 16'b0000001001010001;
    else if (pixel_index == 362 || pixel_index == 383 || pixel_index == 565) oled_data = 16'b0000101001010001;
    else if (pixel_index == 369) oled_data = 16'b0000101001010000;
    else if (pixel_index == 384) oled_data = 16'b0011101011001000;
    else if (pixel_index == 389) oled_data = 16'b0011001001001110;
    else if (pixel_index == 390 || pixel_index == 3267) oled_data = 16'b0011101010001011;
    else if (pixel_index == 391) oled_data = 16'b0011101011001010;
    else if (pixel_index == 393 || pixel_index == 515 || pixel_index == 2474) oled_data = 16'b0101001101000110;
    else if (pixel_index == 394 || pixel_index == 421 || pixel_index == 2184 || pixel_index == 2677) oled_data = 16'b0101001101000100;
    else if (pixel_index == 396 || pixel_index == 1485) oled_data = 16'b0100101101000011;
    else if (pixel_index == 397 || pixel_index == 422 || pixel_index == 517 || pixel_index == 1294 || pixel_index == 1388 || pixel_index == 3515) oled_data = 16'b0100101100000101;
    else if (pixel_index == 399 || pixel_index == 4464 || pixel_index == 4609) oled_data = 16'b0100001011001101;
    else if (pixel_index == 404) oled_data = 16'b0001101001010011;
    else if (pixel_index == 405) oled_data = 16'b0001001001010101;
    else if (pixel_index == 406 || pixel_index == 501) oled_data = 16'b0001101010010101;
    else if (pixel_index == 408 || pixel_index == 503 || pixel_index == 602) oled_data = 16'b0000001001010100;
    else if (pixel_index == 409 || pixel_index == 426 || pixel_index == 525 || pixel_index == 558 || pixel_index == 568 || pixel_index == 668 || pixel_index == 753) oled_data = 16'b0000101001010100;
    else if (pixel_index == 411 || pixel_index == 692) oled_data = 16'b0010001011010100;
    else if (pixel_index == 412) oled_data = 16'b0011001101010100;
    else if (pixel_index == 413) oled_data = 16'b0011101110010001;
    else if (pixel_index == 414) oled_data = 16'b0100001101001111;
    else if (((pixel_index >= 415) && (pixel_index <= 416)) || pixel_index == 927 || pixel_index == 2484) oled_data = 16'b0011101110001100;
    else if (pixel_index == 417) oled_data = 16'b0011101101001101;
    else if (pixel_index == 418) oled_data = 16'b0011101101001010;
    else if (pixel_index == 419 || pixel_index == 1199) oled_data = 16'b0100101110001000;
    else if (pixel_index == 420 || pixel_index == 1198 || pixel_index == 1407 || pixel_index == 2287 || pixel_index == 2572) oled_data = 16'b0101001110000111;
    else if (pixel_index == 425 || pixel_index == 547) oled_data = 16'b0001101010010001;
    else if (pixel_index == 427 || pixel_index == 555 || pixel_index == 746 || pixel_index == 848 || pixel_index == 852) oled_data = 16'b0000001010010100;
    else if (pixel_index == 428) oled_data = 16'b0000101011010010;
    else if (pixel_index == 429) oled_data = 16'b0000001000010100;
    else if (pixel_index == 433 || pixel_index == 534) oled_data = 16'b1001110110101101;
    else if (pixel_index == 434 || pixel_index == 726) oled_data = 16'b0111110101100101;
    else if (pixel_index == 435) oled_data = 16'b0111110101100111;
    else if (pixel_index == 436) oled_data = 16'b0110110100101010;
    else if (pixel_index == 437) oled_data = 16'b0110010010110010;
    else if (pixel_index == 438 || pixel_index == 2036 || pixel_index == 2658) oled_data = 16'b0111010100110010;
    else if (pixel_index == 439 || pixel_index == 1832) oled_data = 16'b1000110101101110;
    else if (pixel_index == 440 || pixel_index == 1737) oled_data = 16'b1000110100101010;
    else if (pixel_index == 441 || pixel_index == 1859 || pixel_index == 1994 || pixel_index == 2171 || pixel_index == 2285) oled_data = 16'b0111010000000100;
    else if (pixel_index == 442 || pixel_index == 1279 || pixel_index == 1508) oled_data = 16'b0110110000000111;
    else if (pixel_index == 443) oled_data = 16'b0110001110001001;
    else if (pixel_index == 444 || pixel_index == 490) oled_data = 16'b0100101100001000;
    else if (pixel_index == 445) oled_data = 16'b0100001011000111;
    else if (pixel_index == 446) oled_data = 16'b0100001100001011;
    else if (pixel_index == 447 || pixel_index == 578 || pixel_index == 688 || pixel_index == 827) oled_data = 16'b0100101100001100;
    else if (pixel_index == 448) oled_data = 16'b0011101011001110;
    else if (pixel_index == 449) oled_data = 16'b0011101100010000;
    else if (pixel_index == 453 || pixel_index == 460 || pixel_index == 463 || pixel_index == 477 || pixel_index == 553 || ((pixel_index >= 556) && (pixel_index <= 557)) || pixel_index == 572 || pixel_index == 654 || pixel_index == 664 || pixel_index == 669) oled_data = 16'b0000101001010011;
    else if (pixel_index == 456) oled_data = 16'b0000001001010000;
    else if (pixel_index == 464 || pixel_index == 554 || pixel_index == 647 || pixel_index == 652) oled_data = 16'b0000001001010011;
    else if (pixel_index == 474 || (pixel_index >= 573) && (pixel_index <= 574)) oled_data = 16'b0001001001010011;
    else if (pixel_index == 483) oled_data = 16'b0100001100001111;
    else if (pixel_index == 484 || pixel_index == 593) oled_data = 16'b0011001011010000;
    else if (pixel_index == 487) oled_data = 16'b0011101101010000;
    else if (pixel_index == 488) oled_data = 16'b0011101100001111;
    else if (pixel_index == 491 || pixel_index == 590 || pixel_index == 1016) oled_data = 16'b0100101101001000;
    else if (pixel_index == 492 || pixel_index == 518) oled_data = 16'b0100101101000101;
    else if (pixel_index == 493 || pixel_index == 999) oled_data = 16'b0011101100000110;
    else if (pixel_index == 494 || pixel_index == 1015 || pixel_index == 1100 || pixel_index == 1936) oled_data = 16'b0100001100000110;
    else if (pixel_index == 495 || pixel_index == 3037) oled_data = 16'b0100101100001011;
    else if (pixel_index == 497) oled_data = 16'b0010001010001111;
    else if (pixel_index == 500 || pixel_index == 549 || pixel_index == 659) oled_data = 16'b0001001010010010;
    else if (pixel_index == 502 || pixel_index == 651) oled_data = 16'b0000101001010101;
    else if (pixel_index == 504 || pixel_index == 601 || pixel_index == 648 || pixel_index == 650 || pixel_index == 655 || pixel_index == 854) oled_data = 16'b0000101010010100;
    else if (pixel_index == 505 || pixel_index == 604 || pixel_index == 697 || pixel_index == 764 || ((pixel_index >= 766) && (pixel_index <= 767)) || pixel_index == 781 || pixel_index == 844 || pixel_index == 858 || ((pixel_index >= 953) && (pixel_index <= 954)) || pixel_index == 958 || pixel_index == 960) oled_data = 16'b0001001011010101;
    else if (pixel_index == 506 || pixel_index == 742 || pixel_index == 744 || pixel_index == 756 || pixel_index == 863) oled_data = 16'b0000101011010100;
    else if (pixel_index == 507 || pixel_index == 561 || pixel_index == 569 || ((pixel_index >= 670) && (pixel_index <= 671)) || pixel_index == 741 || pixel_index == 755 || pixel_index == 760 || pixel_index == 762 || pixel_index == 765) oled_data = 16'b0001001010010100;
    else if (pixel_index == 508 || pixel_index == 843 || pixel_index == 947) oled_data = 16'b0001101100010101;
    else if (pixel_index == 509 || (pixel_index >= 594) && (pixel_index <= 595)) oled_data = 16'b0010001011010010;
    else if (pixel_index == 510) oled_data = 16'b0010001011010000;
    else if (pixel_index == 511 || pixel_index == 608) oled_data = 16'b0010001011001110;
    else if (pixel_index == 512) oled_data = 16'b0001101010001101;
    else if (pixel_index == 513) oled_data = 16'b0010001011001101;
    else if (pixel_index == 514) oled_data = 16'b0011101100001001;
    else if (pixel_index == 516 || pixel_index == 1387 || pixel_index == 1493 || pixel_index == 1672) oled_data = 16'b0101001101000111;
    else if (pixel_index == 520) oled_data = 16'b0010101010001000;
    else if (pixel_index == 522 || pixel_index == 548 || pixel_index == 644) oled_data = 16'b0001101011010001;
    else if (pixel_index == 523 || pixel_index == 700 || pixel_index == 743 || pixel_index == 763 || pixel_index == 859 || ((pixel_index >= 861) && (pixel_index <= 862)) || pixel_index == 956) oled_data = 16'b0001001011010100;
    else if (pixel_index == 524 || pixel_index == 596 || pixel_index == 690) oled_data = 16'b0010001011010011;
    else if (pixel_index == 526 || pixel_index == 993 || pixel_index == 1237) oled_data = 16'b0010001101010101;
    else if (pixel_index == 528 || pixel_index == 675) oled_data = 16'b0100101110001111;
    else if (pixel_index == 529) oled_data = 16'b0111110100101011;
    else if (pixel_index == 530) oled_data = 16'b1000010110101010;
    else if (pixel_index == 531 || pixel_index == 1299) oled_data = 16'b1000010101100101;
    else if (pixel_index == 532) oled_data = 16'b0111010101100111;
    else if (pixel_index == 533 || pixel_index == 1638 || pixel_index == 1848 || pixel_index == 2052 || pixel_index == 2629 || pixel_index == 3065 || pixel_index == 3095) oled_data = 16'b1000010011101100;
    else if (pixel_index == 535) oled_data = 16'b1000010101101001;
    else if (pixel_index == 536 || pixel_index == 2896) oled_data = 16'b0111010011100110;
    else if (pixel_index == 537) oled_data = 16'b0110101111000010;
    else if (pixel_index == 538 || pixel_index == 1412 || pixel_index == 1860 || pixel_index == 3152) oled_data = 16'b0111110000000110;
    else if (pixel_index == 539) oled_data = 16'b0110001110000111;
    else if (pixel_index == 541 || pixel_index == 2580) oled_data = 16'b0011101011000101;
    else if (pixel_index == 542 || pixel_index == 3036) oled_data = 16'b0100101001000111;
    else if (pixel_index == 543) oled_data = 16'b0011101010000110;
    else if (pixel_index == 544 || pixel_index == 641) oled_data = 16'b0011001011001010;
    else if (pixel_index == 545 || pixel_index == 704 || pixel_index == 2977) oled_data = 16'b0011001100001100;
    else if (pixel_index == 546) oled_data = 16'b0010101011001111;
    else if (pixel_index == 559 || pixel_index == 649) oled_data = 16'b0000001001010101;
    else if (pixel_index == 560 || pixel_index == 567 || pixel_index == 646 || pixel_index == 660 || ((pixel_index >= 662) && (pixel_index <= 663)) || pixel_index == 665 || pixel_index == 751 || pixel_index == 761) oled_data = 16'b0000101010010011;
    else if (pixel_index == 562 || pixel_index == 570 || pixel_index == 658 || ((pixel_index >= 666) && (pixel_index <= 667)) || pixel_index == 759) oled_data = 16'b0001001010010011;
    else if (pixel_index == 576) oled_data = 16'b0100001100010000;
    else if (pixel_index == 577 || pixel_index == 5164 || pixel_index == 5167) oled_data = 16'b0100101100001111;
    else if (pixel_index == 579 || pixel_index == 586 || pixel_index == 686 || pixel_index == 1976 || pixel_index == 5264) oled_data = 16'b0100101101001110;
    else if (pixel_index == 584 || pixel_index == 1426) oled_data = 16'b0011101101010001;
    else if (pixel_index == 587 || pixel_index == 3898) oled_data = 16'b0100101110001101;
    else if (pixel_index == 588 || pixel_index == 3897) oled_data = 16'b0100001101001101;
    else if (pixel_index == 591 || pixel_index == 923) oled_data = 16'b0101001100001000;
    else if (pixel_index == 597 || pixel_index == 693 || pixel_index == 842) oled_data = 16'b0001101100010100;
    else if (pixel_index == 598 || pixel_index == 774 || pixel_index == 788 || pixel_index == 882 || pixel_index == 891 || pixel_index == 985 || pixel_index == 1070 || pixel_index == 1088 || pixel_index == 1145 || pixel_index == 1148) oled_data = 16'b0001001100010110;
    else if (pixel_index == 599 || pixel_index == 789 || pixel_index == 876 || pixel_index == 881 || pixel_index == 890 || pixel_index == 984 || pixel_index == 1051) oled_data = 16'b0000101011010110;
    else if (pixel_index == 600 || pixel_index == 745 || pixel_index == 748 || pixel_index == 957) oled_data = 16'b0000101010010101;
    else if (pixel_index == 603 || pixel_index == 835 || pixel_index == 855 || pixel_index == 864) oled_data = 16'b0001001010010101;
    else if (pixel_index == 605 || pixel_index == 679 || pixel_index == 691) oled_data = 16'b0001101011010011;
    else if (pixel_index == 607) oled_data = 16'b0001101010010000;
    else if (pixel_index == 609 || pixel_index == 714) oled_data = 16'b0011001011001001;
    else if (pixel_index == 610) oled_data = 16'b0010001001000100;
    else if (pixel_index == 611) oled_data = 16'b0010101001000001;
    else if (pixel_index == 612) oled_data = 16'b0010101011000011;
    else if (pixel_index == 614 || pixel_index == 809 || pixel_index == 1486 || pixel_index == 1745) oled_data = 16'b0011101011000011;
    else if (pixel_index == 615 || pixel_index == 1581 || pixel_index == 1680 || pixel_index == 2179) oled_data = 16'b0011101100000100;
    else if (pixel_index == 617) oled_data = 16'b0011101011000111;
    else if (pixel_index == 618) oled_data = 16'b0010101101001110;
    else if (pixel_index == 619 || pixel_index == 894) oled_data = 16'b0011101111010100;
    else if (pixel_index == 620 || pixel_index == 1633) oled_data = 16'b0100001111010100;
    else if (pixel_index == 621) oled_data = 16'b0100110001010010;
    else if (pixel_index == 622 || pixel_index == 2115 || pixel_index == 2212 || pixel_index == 2563) oled_data = 16'b0110010010110101;
    else if (pixel_index == 623) oled_data = 16'b1000110110110011;
    else if (pixel_index == 624) oled_data = 16'b1000110110101101;
    else if (pixel_index == 625 || pixel_index == 913) oled_data = 16'b1001111000101011;
    else if (pixel_index == 626 || pixel_index == 816) oled_data = 16'b1001010111101100;
    else if (pixel_index == 627) oled_data = 16'b0111010101100100;
    else if (pixel_index == 628 || pixel_index == 820 || pixel_index == 2995) oled_data = 16'b1000010101100100;
    else if (pixel_index == 629) oled_data = 16'b1000110100100100;
    else if (pixel_index == 630) oled_data = 16'b1001010110100111;
    else if (pixel_index == 631 || pixel_index == 917 || pixel_index == 2521 || pixel_index == 2709) oled_data = 16'b1001010101100110;
    else if (pixel_index == 632 || pixel_index == 1592 || pixel_index == 2618 || pixel_index == 3092) oled_data = 16'b1000110100100110;
    else if (pixel_index == 633 || pixel_index == 1301 || pixel_index == 1574 || pixel_index == 1655 || pixel_index == 1978 || pixel_index == 2766) oled_data = 16'b0110110000000110;
    else if (pixel_index == 634 || pixel_index == 1315 || pixel_index == 1509) oled_data = 16'b0110110001001000;
    else if (pixel_index == 635 || pixel_index == 2033) oled_data = 16'b0110001111001000;
    else if (pixel_index == 636 || pixel_index == 2208) oled_data = 16'b0100101101001010;
    else if (pixel_index == 637) oled_data = 16'b0101001100001011;
    else if (pixel_index == 639 || pixel_index == 709 || pixel_index == 824) oled_data = 16'b0011101011000110;
    else if (pixel_index == 642) oled_data = 16'b0001101010001100;
    else if (pixel_index == 643) oled_data = 16'b0001101010001110;
    else if (pixel_index == 656) oled_data = 16'b0001001011010011;
    else if (pixel_index == 657) oled_data = 16'b0001101010010100;
    else if (pixel_index == 661 || pixel_index == 757) oled_data = 16'b0000101011010011;
    else if (pixel_index == 672) oled_data = 16'b0100001101010011;
    else if (pixel_index == 673) oled_data = 16'b0100101101010100;
    else if (pixel_index == 674) oled_data = 16'b0100001100010001;
    else if (pixel_index == 676 || pixel_index == 1177) oled_data = 16'b0100001110010001;
    else if (pixel_index == 677) oled_data = 16'b0011101100010100;
    else if (pixel_index == 678) oled_data = 16'b0010001011010101;
    else if (pixel_index == 680) oled_data = 16'b0010101100010011;
    else if (pixel_index == 681) oled_data = 16'b0011001101010101;
    else if (pixel_index == 682) oled_data = 16'b0100001101010010;
    else if (pixel_index == 683) oled_data = 16'b0100101110010011;
    else if (pixel_index == 684) oled_data = 16'b0011101101010100;
    else if (pixel_index == 687 || pixel_index == 802 || pixel_index == 1386) oled_data = 16'b0101001101001010;
    else if (((pixel_index >= 694) && (pixel_index <= 695)) || pixel_index == 868) oled_data = 16'b0001001011010110;
    else if (pixel_index == 696 || ((pixel_index >= 776) && (pixel_index <= 777)) || pixel_index == 790 || pixel_index == 873 || pixel_index == 959) oled_data = 16'b0000101011010101;
    else if (pixel_index == 698) oled_data = 16'b0000101100010100;
    else if (pixel_index == 699 || pixel_index == 851 || pixel_index == 865 || pixel_index == 952) oled_data = 16'b0000001011010101;
    else if (pixel_index == 701) oled_data = 16'b0010001100010011;
    else if (pixel_index == 702) oled_data = 16'b0010001100010010;
    else if (pixel_index == 703 || pixel_index == 3844) oled_data = 16'b0010001100001111;
    else if (pixel_index == 705 || pixel_index == 1400 || pixel_index == 1880) oled_data = 16'b0100001100001000;
    else if (pixel_index == 706) oled_data = 16'b0011101100000011;
    else if (pixel_index == 707) oled_data = 16'b0011001011000010;
    else if (pixel_index == 708 || pixel_index == 713) oled_data = 16'b0011101100000101;
    else if (pixel_index == 710) oled_data = 16'b0011001011000101;
    else if (pixel_index == 712 || pixel_index == 1651 || pixel_index == 2176 || pixel_index == 2378) oled_data = 16'b0100101101000100;
    else if (pixel_index == 715) oled_data = 16'b0100101111010000;
    else if (pixel_index == 716) oled_data = 16'b0101010000010000;
    else if (pixel_index == 717 || pixel_index == 1944 || pixel_index == 2037) oled_data = 16'b0110110011110001;
    else if (pixel_index == 718) oled_data = 16'b1001010111110010;
    else if (pixel_index == 719 || pixel_index == 3281) oled_data = 16'b1010111000101111;
    else if (pixel_index == 720) oled_data = 16'b1010011001101011;
    else if (pixel_index == 721 || pixel_index == 818) oled_data = 16'b1001010111101010;
    else if (pixel_index == 722) oled_data = 16'b1010010111101011;
    else if (pixel_index == 723) oled_data = 16'b0111010100100101;
    else if (pixel_index == 724 || pixel_index == 1204) oled_data = 16'b1000110101100101;
    else if (pixel_index == 725) oled_data = 16'b1000110101100100;
    else if (pixel_index == 727 || pixel_index == 1109) oled_data = 16'b0111010011100101;
    else if (pixel_index == 728 || pixel_index == 1476 || pixel_index == 1507 || pixel_index == 1560 || pixel_index == 2269 || pixel_index == 2670) oled_data = 16'b0110110000000101;
    else if (pixel_index == 729 || pixel_index == 1576 || pixel_index == 2483) oled_data = 16'b0100001101000110;
    else if (pixel_index == 730 || pixel_index == 2112 || pixel_index == 3650) oled_data = 16'b0100101101001001;
    else if (pixel_index == 731 || pixel_index == 2819 || pixel_index == 3325) oled_data = 16'b0110001111001010;
    else if (pixel_index == 732) oled_data = 16'b0110110001001010;
    else if (pixel_index == 733) oled_data = 16'b0110110000001100;
    else if (pixel_index == 734 || pixel_index == 1281) oled_data = 16'b0110110001001110;
    else if (pixel_index == 735 || pixel_index == 933 || pixel_index == 2799) oled_data = 16'b0111010001001011;
    else if (pixel_index == 736 || pixel_index == 1380) oled_data = 16'b0110101111001010;
    else if (pixel_index == 737 || pixel_index == 1191) oled_data = 16'b0101001110001101;
    else if (pixel_index == 738) oled_data = 16'b0011001100010000;
    else if (pixel_index == 739) oled_data = 16'b0010001011010001;
    else if (pixel_index == 740 || pixel_index == 786 || pixel_index == 836) oled_data = 16'b0001101011010100;
    else if (pixel_index == 747 || pixel_index == 749 || pixel_index == 849 || pixel_index == 853) oled_data = 16'b0000001010010101;
    else if (pixel_index == 750 || pixel_index == 758) oled_data = 16'b0000001010010011;
    else if (pixel_index == 752) oled_data = 16'b0000101010010010;
    else if (pixel_index == 754) oled_data = 16'b0000101001010110;
    else if (pixel_index == 768) oled_data = 16'b0010101011010110;
    else if (pixel_index == 769) oled_data = 16'b0011001011010100;
    else if (pixel_index == 770) oled_data = 16'b0011001100010100;
    else if (pixel_index == 771) oled_data = 16'b0100001110010011;
    else if (pixel_index == 772 || pixel_index == 930 || pixel_index == 2498) oled_data = 16'b0011101110010011;
    else if (pixel_index == 773 || pixel_index == 1619) oled_data = 16'b0010101110010110;
    else if (pixel_index == 775 || pixel_index == 874 || pixel_index == 949 || pixel_index == 987 || pixel_index == 1084) oled_data = 16'b0000101100010111;
    else if (pixel_index == 778) oled_data = 16'b0010001100010110;
    else if (pixel_index == 779) oled_data = 16'b0010101100010101;
    else if (pixel_index == 780 || pixel_index == 1047) oled_data = 16'b0001101100010110;
    else if (pixel_index == 782) oled_data = 16'b0011001100010011;
    else if (pixel_index == 783) oled_data = 16'b0011101100010010;
    else if (pixel_index == 784) oled_data = 16'b0100101011010011;
    else if (pixel_index == 785) oled_data = 16'b0011001011010101;
    else if (pixel_index == 787 || pixel_index == 834) oled_data = 16'b0001001100010100;
    else if (pixel_index == 791 || pixel_index == 846 || pixel_index == 883 || pixel_index == 888) oled_data = 16'b0000101100010101;
    else if (pixel_index == 792 || (pixel_index >= 794) && (pixel_index <= 795)) oled_data = 16'b0000101101010101;
    else if (pixel_index == 793 || pixel_index == 872 || pixel_index == 885 || pixel_index == 889 || pixel_index == 972 || pixel_index == 1052 || pixel_index == 1054 || pixel_index == 1238) oled_data = 16'b0000001100010110;
    else if (pixel_index == 796 || pixel_index == 982 || pixel_index == 1048) oled_data = 16'b0001001101010101;
    else if (pixel_index == 797) oled_data = 16'b0010001110010011;
    else if (pixel_index == 798) oled_data = 16'b0011001110010010;
    else if (pixel_index == 799) oled_data = 16'b0100001110001111;
    else if (pixel_index == 800 || pixel_index == 3269) oled_data = 16'b0101101110001100;
    else if (pixel_index == 801) oled_data = 16'b0110101111001100;
    else if (pixel_index == 804) oled_data = 16'b0100101111001010;
    else if (pixel_index == 805 || pixel_index == 2373 || pixel_index == 2566 || pixel_index == 3747) oled_data = 16'b0101001111001001;
    else if (pixel_index == 807 || pixel_index == 2374) oled_data = 16'b0100101110000101;
    else if (pixel_index == 808 || pixel_index == 2079) oled_data = 16'b0100101100000010;
    else if (pixel_index == 810) oled_data = 16'b0010001001000101;
    else if (pixel_index == 812 || pixel_index == 1023) oled_data = 16'b0101001111001100;
    else if (pixel_index == 813) oled_data = 16'b0110110011101110;
    else if (pixel_index == 814) oled_data = 16'b1000110111110000;
    else if (pixel_index == 815) oled_data = 16'b1001110111101111;
    else if (pixel_index == 817) oled_data = 16'b1000110110101001;
    else if (pixel_index == 819) oled_data = 16'b0110110100100011;
    else if (pixel_index == 821 || pixel_index == 3091) oled_data = 16'b1000110110100101;
    else if (pixel_index == 822 || pixel_index == 2524 || pixel_index == 2620) oled_data = 16'b1000010100100101;
    else if (pixel_index == 823 || pixel_index == 1649 || pixel_index == 2470) oled_data = 16'b0101001111000101;
    else if (pixel_index == 825 || pixel_index == 1210) oled_data = 16'b0001001001001010;
    else if (pixel_index == 828 || pixel_index == 1289) oled_data = 16'b0101101110001011;
    else if (pixel_index == 829 || pixel_index == 1977) oled_data = 16'b0101001101001000;
    else if (pixel_index == 830) oled_data = 16'b0100101110001001;
    else if (pixel_index == 831) oled_data = 16'b0101101111001100;
    else if (pixel_index == 832) oled_data = 16'b0101101110001110;
    else if (pixel_index == 838) oled_data = 16'b0001101011010010;
    else if (pixel_index == 839) oled_data = 16'b0010001101010100;
    else if (pixel_index == 840) oled_data = 16'b0010101101010100;
    else if (pixel_index == 841) oled_data = 16'b0010001100010100;
    else if (pixel_index == 845 || pixel_index == 964) oled_data = 16'b0000001100010101;
    else if (pixel_index == 847 || pixel_index == 860 || pixel_index == 955) oled_data = 16'b0001001100010101;
    else if (pixel_index == 850) oled_data = 16'b0000001010010110;
    else if (((pixel_index >= 856) && (pixel_index <= 857)) || pixel_index == 867) oled_data = 16'b0001001010010110;
    else if (pixel_index == 866 || pixel_index == 948 || ((pixel_index >= 965) && (pixel_index <= 966)) || pixel_index == 983 || pixel_index == 986 || pixel_index == 1050 || pixel_index == 1146) oled_data = 16'b0000101100010110;
    else if (((pixel_index >= 869) && (pixel_index <= 870)) || pixel_index == 1058 || pixel_index == 1063 || pixel_index == 1066 || pixel_index == 1155 || pixel_index == 1172 || pixel_index == 1244) oled_data = 16'b0001001110010111;
    else if (pixel_index == 871 || pixel_index == 1046 || pixel_index == 1089 || pixel_index == 1334) oled_data = 16'b0001101101010111;
    else if (pixel_index == 875) oled_data = 16'b0000001010010111;
    else if (pixel_index == 877 || pixel_index == 1069 || pixel_index == 1255) oled_data = 16'b0000001101010111;
    else if (pixel_index == 878 || pixel_index == 981 || pixel_index == 1082 || pixel_index == 1158) oled_data = 16'b0001001110010110;
    else if (pixel_index == 879 || pixel_index == 1062 || pixel_index == 1072 || pixel_index == 1142 || pixel_index == 1147 || pixel_index == 1149 || pixel_index == 1151 || pixel_index == 1248 || pixel_index == 1335) oled_data = 16'b0001001101010111;
    else if (pixel_index == 880 || pixel_index == 950 || pixel_index == 968) oled_data = 16'b0001001100010111;
    else if (pixel_index == 884 || pixel_index == 961 || pixel_index == 971 || pixel_index == 1086 || pixel_index == 1159) oled_data = 16'b0000101101010110;
    else if (pixel_index == 886) oled_data = 16'b0000001011010100;
    else if (pixel_index == 887) oled_data = 16'b0000001101010101;
    else if (pixel_index == 892 || pixel_index == 980 || pixel_index == 1071 || pixel_index == 1081 || ((pixel_index >= 1143) && (pixel_index <= 1144)) || pixel_index == 1150) oled_data = 16'b0001001101010110;
    else if (pixel_index == 893) oled_data = 16'b0010001110010101;
    else if (pixel_index == 895 || pixel_index == 943 || pixel_index == 1287 || pixel_index == 2239) oled_data = 16'b0110110001010000;
    else if (pixel_index == 896 || pixel_index == 2069) oled_data = 16'b0111010000001111;
    else if (pixel_index == 897) oled_data = 16'b0101101110010001;
    else if (pixel_index == 898 || pixel_index == 5080) oled_data = 16'b0101101111010011;
    else if (pixel_index == 899 || pixel_index == 2240 || pixel_index == 3126) oled_data = 16'b0111010011110001;
    else if (pixel_index == 900) oled_data = 16'b0110010011101100;
    else if (pixel_index == 901) oled_data = 16'b0110010001001010;
    else if (pixel_index == 902 || pixel_index == 1422 || pixel_index == 1693 || pixel_index == 2576) oled_data = 16'b0101110000001000;
    else if (pixel_index == 903) oled_data = 16'b0011101101000100;
    else if (pixel_index == 904 || pixel_index == 1391) oled_data = 16'b0010101010000001;
    else if (pixel_index == 905) oled_data = 16'b0001101001000001;
    else if (pixel_index == 906) oled_data = 16'b0010001001000010;
    else if (pixel_index == 907) oled_data = 16'b0011101001000100;
    else if (pixel_index == 910) oled_data = 16'b0111110110101100;
    else if (pixel_index == 911) oled_data = 16'b0101110010101001;
    else if (pixel_index == 912) oled_data = 16'b1000111000101011;
    else if (pixel_index == 914) oled_data = 16'b1001010101101010;
    else if (pixel_index == 915) oled_data = 16'b0110110101100001;
    else if (pixel_index == 916) oled_data = 16'b0111010101100011;
    else if (pixel_index == 918 || pixel_index == 2088 || pixel_index == 2092) oled_data = 16'b0110001110000100;
    else if (pixel_index == 919 || pixel_index == 1019 || pixel_index == 1113) oled_data = 16'b0010001001000110;
    else if (pixel_index == 920) oled_data = 16'b0010101011000111;
    else if (pixel_index == 921) oled_data = 16'b0100001110001011;
    else if (pixel_index == 922) oled_data = 16'b0110010000001101;
    else if (pixel_index == 925 || pixel_index == 1584 || pixel_index == 3226) oled_data = 16'b0010101001000011;
    else if (pixel_index == 928) oled_data = 16'b0100001111001111;
    else if (pixel_index == 929 || pixel_index == 3899) oled_data = 16'b0100001111010001;
    else if (pixel_index == 931 || pixel_index == 2062 || pixel_index == 2661) oled_data = 16'b0101010001010010;
    else if (pixel_index == 932 || pixel_index == 996 || pixel_index == 1288 || pixel_index == 2535) oled_data = 16'b0111010001001110;
    else if (pixel_index == 934 || pixel_index == 1647 || pixel_index == 1675 || pixel_index == 2630) oled_data = 16'b0111010001001010;
    else if (pixel_index == 935) oled_data = 16'b1010010101101111;
    else if (pixel_index == 936) oled_data = 16'b1010110101101110;
    else if (pixel_index == 937) oled_data = 16'b1001010011101110;
    else if (pixel_index == 938 || pixel_index == 2908) oled_data = 16'b1001010101101110;
    else if (pixel_index == 939) oled_data = 16'b1000010011110000;
    else if (pixel_index == 941 || pixel_index == 1519 || pixel_index == 2559 || pixel_index == 4899) oled_data = 16'b0111010010110000;
    else if (pixel_index == 942 || pixel_index == 1286 || pixel_index == 2553) oled_data = 16'b0110010000010001;
    else if (pixel_index == 944 || pixel_index == 2883) oled_data = 16'b0100101110010010;
    else if (pixel_index == 945) oled_data = 16'b0011001101010010;
    else if (pixel_index == 946) oled_data = 16'b0010001101010011;
    else if (pixel_index == 951) oled_data = 16'b0000101011010111;
    else if (pixel_index == 962 || ((pixel_index >= 975) && (pixel_index <= 976)) || pixel_index == 1083 || pixel_index == 1154 || pixel_index == 1165 || pixel_index == 1239 || pixel_index == 1246) oled_data = 16'b0000101101010111;
    else if (pixel_index == 963 || pixel_index == 969 || pixel_index == 988 || (pixel_index >= 1079) && (pixel_index <= 1080)) oled_data = 16'b0000001100010111;
    else if (pixel_index == 967 || pixel_index == 1057 || pixel_index == 1245 || ((pixel_index >= 1249) && (pixel_index <= 1250)) || pixel_index == 1339 || pixel_index == 1347 || ((pixel_index >= 1435) && (pixel_index <= 1436)) || ((pixel_index >= 1438) && (pixel_index <= 1439)) || pixel_index == 1444) oled_data = 16'b0001001101011000;
    else if (pixel_index == 970) oled_data = 16'b0000001101010110;
    else if (pixel_index == 973 || pixel_index == 977 || pixel_index == 979 || pixel_index == 989 || pixel_index == 1074 || pixel_index == 1076 || pixel_index == 1160 || pixel_index == 1163 || pixel_index == 1240 || pixel_index == 1242) oled_data = 16'b0000101101011000;
    else if (pixel_index == 974 || pixel_index == 1056 || pixel_index == 1064) oled_data = 16'b0000101100011000;
    else if (pixel_index == 978 || pixel_index == 1167 || pixel_index == 1254 || pixel_index == 1346) oled_data = 16'b0000101110011000;
    else if (pixel_index == 990 || pixel_index == 1184 || pixel_index == 1243 || pixel_index == 1247 || pixel_index == 1333) oled_data = 16'b0001101101010110;
    else if (pixel_index == 991 || pixel_index == 1179) oled_data = 16'b0100101111010001;
    else if (pixel_index == 992) oled_data = 16'b0011001110010011;
    else if (pixel_index == 994) oled_data = 16'b0011101111010111;
    else if (pixel_index == 995) oled_data = 16'b0110010001010100;
    else if (pixel_index == 997 || pixel_index == 1742 || pixel_index == 2718 || pixel_index == 2860 || pixel_index == 2865) oled_data = 16'b0111010010101100;
    else if (pixel_index == 998 || pixel_index == 1094 || pixel_index == 1938) oled_data = 16'b0110010000001010;
    else if (pixel_index == 1000) oled_data = 16'b0010101001000100;
    else if (pixel_index == 1002 || pixel_index == 1786 || pixel_index == 2279) oled_data = 16'b0101101110000100;
    else if (pixel_index == 1003 || pixel_index == 1985 || pixel_index == 2080) oled_data = 16'b0100001011000010;
    else if (pixel_index == 1006) oled_data = 16'b1001010111101011;
    else if (pixel_index == 1007) oled_data = 16'b0101110011101000;
    else if (pixel_index == 1008) oled_data = 16'b1000010101101011;
    else if (pixel_index == 1009) oled_data = 16'b1010111001101110;
    else if (pixel_index == 1010 || pixel_index == 1214) oled_data = 16'b1010011000101100;
    else if (pixel_index == 1011) oled_data = 16'b1000110111100010;
    else if (pixel_index == 1012) oled_data = 16'b0111010011100011;
    else if (pixel_index == 1013 || pixel_index == 1475 || pixel_index == 1568 || pixel_index == 1757 || pixel_index == 1867 || pixel_index == 1958 || pixel_index == 2612) oled_data = 16'b1000010001000101;
    else if (pixel_index == 1014) oled_data = 16'b0101110000000100;
    else if (pixel_index == 1018) oled_data = 16'b0011101001000111;
    else if (pixel_index == 1020) oled_data = 16'b0010001010000101;
    else if (pixel_index == 1021 || pixel_index == 2940) oled_data = 16'b0011001001000101;
    else if (pixel_index == 1022 || pixel_index == 3129) oled_data = 16'b0011001010000101;
    else if (pixel_index == 1024 || pixel_index == 1773 || pixel_index == 2467 || pixel_index == 3518) oled_data = 16'b0111010010101110;
    else if (pixel_index == 1025) oled_data = 16'b1010010110101111;
    else if (pixel_index == 1026) oled_data = 16'b1001110101101111;
    else if (pixel_index == 1027) oled_data = 16'b1001110111101011;
    else if (pixel_index == 1028 || pixel_index == 1032) oled_data = 16'b1010110111101000;
    else if (pixel_index == 1029 || pixel_index == 2428) oled_data = 16'b1000110100100101;
    else if (pixel_index == 1030 || pixel_index == 1125) oled_data = 16'b0111110010100101;
    else if (pixel_index == 1031) oled_data = 16'b1001010100101001;
    else if (pixel_index == 1033 || pixel_index == 1736) oled_data = 16'b1010010110101000;
    else if (pixel_index == 1034) oled_data = 16'b1010010110100111;
    else if (pixel_index == 1035) oled_data = 16'b1001110100100111;
    else if (pixel_index == 1036 || pixel_index == 1123 || pixel_index == 1129 || pixel_index == 2707) oled_data = 16'b1001010100101000;
    else if (pixel_index == 1037 || pixel_index == 1643 || pixel_index == 1896 || pixel_index == 1898 || pixel_index == 2897) oled_data = 16'b1000110100101001;
    else if (pixel_index == 1038 || pixel_index == 1378 || pixel_index == 1868 || pixel_index == 2465 || pixel_index == 2561 || pixel_index == 3000 || pixel_index == 3063 || pixel_index == 4128) oled_data = 16'b0111010000001000;
    else if (pixel_index == 1039 || pixel_index == 1321 || pixel_index == 3157) oled_data = 16'b0110110000001001;
    else if (pixel_index == 1040 || pixel_index == 1270) oled_data = 16'b1000010010101100;
    else if (pixel_index == 1041 || pixel_index == 2144 || (pixel_index >= 3252) && (pixel_index <= 3253)) oled_data = 16'b1000110011101110;
    else if (pixel_index == 1042 || pixel_index == 1922) oled_data = 16'b0111110010110001;
    else if (pixel_index == 1043 || pixel_index == 3903) oled_data = 16'b0100010000010101;
    else if (pixel_index == 1044) oled_data = 16'b0010001100010111;
    else if (pixel_index == 1045) oled_data = 16'b0001101100010111;
    else if (pixel_index == 1049) oled_data = 16'b0001001110010100;
    else if (pixel_index == 1053 || pixel_index == 1055 || pixel_index == 1060) oled_data = 16'b0000001011010110;
    else if (pixel_index == 1059) oled_data = 16'b0000001110010111;
    else if (pixel_index == 1061) oled_data = 16'b0000001011010111;
    else if (pixel_index == 1065 || pixel_index == 1337 || pixel_index == 1341 || (pixel_index >= 1533) && (pixel_index <= 1534)) oled_data = 16'b0001001110011001;
    else if ((pixel_index >= 1067) && (pixel_index <= 1068)) oled_data = 16'b0000101110010110;
    else if (pixel_index == 1073 || pixel_index == 1164 || pixel_index == 1170 || pixel_index == 1173 || pixel_index == 1348) oled_data = 16'b0000101110010111;
    else if (pixel_index == 1075 || pixel_index == 1153 || pixel_index == 1166) oled_data = 16'b0000001101011000;
    else if (pixel_index == 1077 || pixel_index == 1085) oled_data = 16'b0000001100011000;
    else if (pixel_index == 1078) oled_data = 16'b0000001011011000;
    else if (pixel_index == 1087) oled_data = 16'b0011001110010101;
    else if (pixel_index == 1090) oled_data = 16'b0100001110010111;
    else if (pixel_index == 1091 || pixel_index == 4988) oled_data = 16'b0111010000010100;
    else if (pixel_index == 1092 || pixel_index == 2159 || pixel_index == 3098 || pixel_index == 3272) oled_data = 16'b1000010001001111;
    else if (pixel_index == 1093 || pixel_index == 2151 || pixel_index == 2194 || pixel_index == 2464 || pixel_index == 2797 || pixel_index == 4224) oled_data = 16'b0111110010101101;
    else if (pixel_index == 1096) oled_data = 16'b0011001010000011;
    else if (pixel_index == 1097) oled_data = 16'b0101101011000101;
    else if (pixel_index == 1098) oled_data = 16'b0100101010000101;
    else if (pixel_index == 1099) oled_data = 16'b0011001000000100;
    else if (pixel_index == 1101 || pixel_index == 1489) oled_data = 16'b0001101000000011;
    else if (pixel_index == 1102 || pixel_index == 1492 || pixel_index == 2803) oled_data = 16'b1000010011100111;
    else if (pixel_index == 1103 || pixel_index == 1325 || pixel_index == 1885 || pixel_index == 2675) oled_data = 16'b0101110000000110;
    else if (pixel_index == 1104) oled_data = 16'b0111110100101000;
    else if (pixel_index == 1105) oled_data = 16'b1010111010101111;
    else if (pixel_index == 1106) oled_data = 16'b1011111001101101;
    else if (pixel_index == 1107) oled_data = 16'b1001111000100010;
    else if (pixel_index == 1108) oled_data = 16'b0101110001000011;
    else if (pixel_index == 1110 || pixel_index == 1414 || pixel_index == 2811) oled_data = 16'b0111110010100110;
    else if (pixel_index == 1111 || pixel_index == 1377 || pixel_index == 1750) oled_data = 16'b0110001111000111;
    else if (pixel_index == 1112) oled_data = 16'b0011001010001000;
    else if (pixel_index == 1114) oled_data = 16'b0001101000001010;
    else if (pixel_index == 1117) oled_data = 16'b0100101110001010;
    else if (pixel_index == 1118 || pixel_index == 1479 || pixel_index == 2864) oled_data = 16'b0111010010101010;
    else if (pixel_index == 1119) oled_data = 16'b1010111000101100;
    else if (pixel_index == 1120 || pixel_index == 1319 || pixel_index == 2244) oled_data = 16'b1010010101101010;
    else if (pixel_index == 1121) oled_data = 16'b1100011000101010;
    else if (pixel_index == 1122) oled_data = 16'b1011111000101011;
    else if (pixel_index == 1124) oled_data = 16'b1001010011100101;
    else if (pixel_index == 1126 || pixel_index == 1471 || pixel_index == 1567 || pixel_index == 2190) oled_data = 16'b0111010001000101;
    else if (pixel_index == 1127 || pixel_index == 1363 || pixel_index == 1548 || pixel_index == 1950) oled_data = 16'b1001010011101000;
    else if (pixel_index == 1128 || pixel_index == 1130) oled_data = 16'b1001110100101001;
    else if (pixel_index == 1131 || pixel_index == 1362) oled_data = 16'b1001010100100111;
    else if (pixel_index == 1132 || pixel_index == 1499 || pixel_index == 2433 || pixel_index == 2518 || pixel_index == 2522) oled_data = 16'b1001110101100111;
    else if (pixel_index == 1133 || pixel_index == 2336 || pixel_index == 2432 || pixel_index == 2625) oled_data = 16'b1001110101101000;
    else if (pixel_index == 1134 || pixel_index == 1644) oled_data = 16'b1000010011101010;
    else if (pixel_index == 1135 || pixel_index == 2209) oled_data = 16'b0101001110001011;
    else if (pixel_index == 1136 || pixel_index == 3320 || pixel_index == 5991 || pixel_index == 6049 || pixel_index == 6059) oled_data = 16'b0110101110001111;
    else if (pixel_index == 1137) oled_data = 16'b1000110011110000;
    else if (pixel_index == 1138 || pixel_index == 2699 || pixel_index == 2890 || pixel_index == 3270) oled_data = 16'b0111110011110011;
    else if (pixel_index == 1139) oled_data = 16'b0101010000010101;
    else if (pixel_index == 1140) oled_data = 16'b0001101110010110;
    else if (pixel_index == 1141 || pixel_index == 1157) oled_data = 16'b0001001100011000;
    else if (pixel_index == 1152 || pixel_index == 1257) oled_data = 16'b0000001101011001;
    else if (pixel_index == 1156 || pixel_index == 1161) oled_data = 16'b0001001101011001;
    else if (pixel_index == 1162) oled_data = 16'b0000101110011001;
    else if (((pixel_index >= 1168) && (pixel_index <= 1169)) || pixel_index == 1256) oled_data = 16'b0000001110011000;
    else if (pixel_index == 1171 || pixel_index == 1336 || pixel_index == 1340 || pixel_index == 1343) oled_data = 16'b0001101110011000;
    else if (pixel_index == 1174 || pixel_index == 1445) oled_data = 16'b0010001110010111;
    else if (pixel_index == 1175 || pixel_index == 1355 || pixel_index == 1795 || pixel_index == 2786) oled_data = 16'b0011110000010101;
    else if (pixel_index == 1176) oled_data = 16'b0011101111010010;
    else if (pixel_index == 1178) oled_data = 16'b0100101111010010;
    else if (pixel_index == 1180) oled_data = 16'b0101001101010001;
    else if (pixel_index == 1181 || pixel_index == 5078) oled_data = 16'b0101001110010010;
    else if (pixel_index == 1182 || pixel_index == 3902) oled_data = 16'b0011101111010011;
    else if (pixel_index == 1183) oled_data = 16'b0010101111010010;
    else if (pixel_index == 1185 || pixel_index == 1251) oled_data = 16'b0001101110010111;
    else if (pixel_index == 1186) oled_data = 16'b0010001101010110;
    else if (pixel_index == 1187) oled_data = 16'b0011101101010111;
    else if (pixel_index == 1188) oled_data = 16'b0101001110010100;
    else if (pixel_index == 1189 || pixel_index == 2129) oled_data = 16'b0101010000010010;
    else if (pixel_index == 1192 || pixel_index == 2153) oled_data = 16'b1000001111001010;
    else if (pixel_index == 1193 || pixel_index == 2822) oled_data = 16'b0101101101001000;
    else if (pixel_index == 1194) oled_data = 16'b0100001001000110;
    else if (pixel_index == 1195 || pixel_index == 1302) oled_data = 16'b0010101000000011;
    else if (pixel_index == 1196 || pixel_index == 3649) oled_data = 16'b0101001011000011;
    else if (pixel_index == 1197) oled_data = 16'b0100001011000001;
    else if (pixel_index == 1200) oled_data = 16'b0100110000000111;
    else if (pixel_index == 1201 || pixel_index == 1307 || pixel_index == 1480 || pixel_index == 2717) oled_data = 16'b1000010100101100;
    else if (pixel_index == 1203) oled_data = 16'b1001110111100101;
    else if (pixel_index == 1205 || pixel_index == 1491) oled_data = 16'b0111010010100100;
    else if (pixel_index == 1206 || pixel_index == 1588) oled_data = 16'b0100001100000101;
    else if (pixel_index == 1208) oled_data = 16'b0010100111000101;
    else if (pixel_index == 1209) oled_data = 16'b0001100110000111;
    else if (pixel_index == 1211) oled_data = 16'b0011001111010001;
    else if (pixel_index == 1212 || pixel_index == 2020 || pixel_index == 2439 || pixel_index == 3653) oled_data = 16'b0110110011110010;
    else if (pixel_index == 1213) oled_data = 16'b1001010110101110;
    else if (pixel_index == 1215) oled_data = 16'b1100111001101011;
    else if (pixel_index == 1216) oled_data = 16'b1000110101101001;
    else if (pixel_index == 1217) oled_data = 16'b1000010100101001;
    else if (pixel_index == 1218) oled_data = 16'b1011010110101010;
    else if (pixel_index == 1219 || pixel_index == 1273 || pixel_index == 1685 || pixel_index == 2422 || pixel_index == 3158) oled_data = 16'b0111110001001000;
    else if (pixel_index == 1220 || pixel_index == 1648 || pixel_index == 1762) oled_data = 16'b0110010001000101;
    else if (pixel_index == 1221) oled_data = 16'b0111010010100110;
    else if (pixel_index == 1222) oled_data = 16'b1000010011100101;
    else if (pixel_index == 1223) oled_data = 16'b1010110110101011;
    else if (pixel_index == 1224 || pixel_index == 1949) oled_data = 16'b1001110011101011;
    else if (pixel_index == 1225 || pixel_index == 1401 || pixel_index == 1495 || pixel_index == 1741) oled_data = 16'b0111110010101001;
    else if (pixel_index == 1226 || pixel_index == 1230) oled_data = 16'b1010010011101000;
    else if (pixel_index == 1227 || pixel_index == 1370 || pixel_index == 1562 || pixel_index == 1658 || pixel_index == 2610) oled_data = 16'b1000010010100110;
    else if (pixel_index == 1228 || pixel_index == 1456 || pixel_index == 2425 || pixel_index == 2517) oled_data = 16'b1001010011100111;
    else if (pixel_index == 1229 || pixel_index == 2516 || pixel_index == 2617) oled_data = 16'b1000110010100110;
    else if (pixel_index == 1231 || pixel_index == 1947) oled_data = 16'b1000010001001011;
    else if (pixel_index == 1232 || pixel_index == 2210) oled_data = 16'b0101101111001111;
    else if (pixel_index == 1233 || pixel_index == 3996) oled_data = 16'b0100110000010010;
    else if (pixel_index == 1234 || pixel_index == 2222 || pixel_index == 3995) oled_data = 16'b0101010001010011;
    else if (pixel_index == 1235 || pixel_index == 2158) oled_data = 16'b0101110001010100;
    else if (pixel_index == 1236 || pixel_index == 1702 || pixel_index == 2359) oled_data = 16'b0011101111010101;
    else if (pixel_index == 1241) oled_data = 16'b0000101101011001;
    else if (pixel_index == 1252 || pixel_index == 1530) oled_data = 16'b0001001111011000;
    else if (pixel_index == 1253 || pixel_index == 1537 || (pixel_index >= 1627) && (pixel_index <= 1628)) oled_data = 16'b0001001111011001;
    else if ((pixel_index >= 1258) && (pixel_index <= 1259)) oled_data = 16'b0000001110011001;
    else if (pixel_index == 1260 || pixel_index == 1338 || pixel_index == 1345 || pixel_index == 1434 || pixel_index == 1437 || pixel_index == 1535) oled_data = 16'b0001001110011000;
    else if (pixel_index == 1261) oled_data = 16'b0010001110011000;
    else if (pixel_index == 1262 || pixel_index == 1331) oled_data = 16'b0011001111010101;
    else if (pixel_index == 1263 || pixel_index == 1729) oled_data = 16'b0100010000010100;
    else if (pixel_index == 1264 || pixel_index == 2120 || pixel_index == 2663) oled_data = 16'b0101110010110000;
    else if (pixel_index == 1265 || pixel_index == 1694 || pixel_index == 1940 || pixel_index == 2028 || pixel_index == 2510) oled_data = 16'b0110010010101111;
    else if (pixel_index == 1266 || pixel_index == 2026) oled_data = 16'b0101110001001110;
    else if (pixel_index == 1267 || pixel_index == 2861) oled_data = 16'b0110010001001111;
    else if (pixel_index == 1268) oled_data = 16'b0110110001001100;
    else if (pixel_index == 1269 || pixel_index == 1834 || pixel_index == 1837 || pixel_index == 2674 || pixel_index == 2962) oled_data = 16'b0110110010101100;
    else if (pixel_index == 1271 || pixel_index == 1320) oled_data = 16'b1000110011101011;
    else if (pixel_index == 1272 || pixel_index == 1853 || pixel_index == 2054) oled_data = 16'b1000010010101001;
    else if (pixel_index == 1274 || pixel_index == 1876) oled_data = 16'b0111110010100111;
    else if (pixel_index == 1275 || pixel_index == 1755) oled_data = 16'b0111010000000111;
    else if (pixel_index == 1276 || pixel_index == 3056) oled_data = 16'b0110101111000111;
    else if (pixel_index == 1277 || pixel_index == 2702 || pixel_index == 2960 || pixel_index == 3422) oled_data = 16'b0110101111001001;
    else if (pixel_index == 1280 || pixel_index == 3421) oled_data = 16'b0111010000001011;
    else if (pixel_index == 1282 || pixel_index == 2605) oled_data = 16'b0110010000001111;
    else if (pixel_index == 1283 || pixel_index == 1607 || pixel_index == 2024) oled_data = 16'b0110010001010001;
    else if (((pixel_index >= 1284) && (pixel_index <= 1285)) || pixel_index == 2211) oled_data = 16'b0110010000010010;
    else if (pixel_index == 1290) oled_data = 16'b0100101010000111;
    else if (pixel_index == 1291 || pixel_index == 1390 || pixel_index == 3457) oled_data = 16'b0100001010000011;
    else if (pixel_index == 1292) oled_data = 16'b0101001100000011;
    else if (pixel_index == 1293 || pixel_index == 2476) oled_data = 16'b0101001101000101;
    else if (pixel_index == 1295) oled_data = 16'b0011001100000110;
    else if (pixel_index == 1296) oled_data = 16'b0101010001000101;
    else if (pixel_index == 1297) oled_data = 16'b1000110101101010;
    else if (pixel_index == 1298) oled_data = 16'b1011011011101111;
    else if (pixel_index == 1300 || pixel_index == 2436 || pixel_index == 2626 || pixel_index == 2710) oled_data = 16'b1001010101100111;
    else if (pixel_index == 1303) oled_data = 16'b0001000101000001;
    else if (pixel_index == 1304 || pixel_index == 3025) oled_data = 16'b0010000101000011;
    else if (pixel_index == 1305 || pixel_index == 2731) oled_data = 16'b0011001000000101;
    else if (pixel_index == 1308) oled_data = 16'b1010011000101011;
    else if (pixel_index == 1309) oled_data = 16'b1011011000101010;
    else if (pixel_index == 1310) oled_data = 16'b1010010110101010;
    else if (pixel_index == 1311) oled_data = 16'b1011010101101011;
    else if (pixel_index == 1312) oled_data = 16'b1001110100101011;
    else if (pixel_index == 1313 || pixel_index == 1478 || pixel_index == 1846 || pixel_index == 1878) oled_data = 16'b0110110000001000;
    else if (pixel_index == 1314 || pixel_index == 1642 || pixel_index == 2193 || pixel_index == 3159) oled_data = 16'b1000010011101001;
    else if (pixel_index == 1316 || pixel_index == 1371 || ((pixel_index >= 2093) && (pixel_index <= 2094)) || pixel_index == 2772) oled_data = 16'b0110010000000101;
    else if (pixel_index == 1317) oled_data = 16'b0110110001000101;
    else if (pixel_index == 1318 || pixel_index == 1563 || pixel_index == 1659 || pixel_index == 2366) oled_data = 16'b0111110001000101;
    else if (pixel_index == 1322 || pixel_index == 1753) oled_data = 16'b1000110010101001;
    else if (pixel_index == 1323) oled_data = 16'b0111001111000110;
    else if (pixel_index == 1324) oled_data = 16'b0111010001000111;
    else if (pixel_index == 1326) oled_data = 16'b0110110010100111;
    else if (pixel_index == 1327 || pixel_index == 1561 || pixel_index == 2051) oled_data = 16'b1000010010100111;
    else if (pixel_index == 1328 || pixel_index == 1743 || pixel_index == 1932) oled_data = 16'b0110010000001100;
    else if (pixel_index == 1329) oled_data = 16'b0011101111010001;
    else if (pixel_index == 1330) oled_data = 16'b0011001111010010;
    else if (pixel_index == 1332) oled_data = 16'b0011001111010110;
    else if (pixel_index == 1342) oled_data = 16'b0001101101011000;
    else if (pixel_index == 1344) oled_data = 16'b0000101111010111;
    else if (pixel_index == 1349) oled_data = 16'b0000001111011001;
    else if (pixel_index == 1350 || pixel_index == 1441 || pixel_index == 1706) oled_data = 16'b0000101111011010;
    else if (pixel_index == 1351) oled_data = 16'b0000101111011011;
    else if (pixel_index == 1352 || pixel_index == 1622 || pixel_index == 1705 || ((pixel_index >= 1719) && (pixel_index <= 1720)) || pixel_index == 1805 || pixel_index == 1815 || pixel_index == 1817 || pixel_index == 1819 || pixel_index == 1916) oled_data = 16'b0001110000011010;
    else if (pixel_index == 1353 || (pixel_index >= 3911) && (pixel_index <= 3913)) oled_data = 16'b0001101111010110;
    else if (pixel_index == 1354 || pixel_index == 2688) oled_data = 16'b0010110000010100;
    else if (pixel_index == 1356 || pixel_index == 2219 || pixel_index == 2918) oled_data = 16'b0101010010110100;
    else if (pixel_index == 1357 || pixel_index == 2041) oled_data = 16'b0110110011110011;
    else if (pixel_index == 1358 || pixel_index == 1500) oled_data = 16'b1001010100101011;
    else if (pixel_index == 1359 || pixel_index == 2519 || pixel_index == 2528) oled_data = 16'b1010010100100111;
    else if (pixel_index == 1360) oled_data = 16'b1010110101100011;
    else if (pixel_index == 1361) oled_data = 16'b1010110100100110;
    else if (pixel_index == 1364 || pixel_index == 1455 || pixel_index == 1469 || pixel_index == 1547 || pixel_index == 1570) oled_data = 16'b1001110011100110;
    else if (pixel_index == 1365) oled_data = 16'b1010010101100110;
    else if (pixel_index == 1366) oled_data = 16'b1010110011100111;
    else if (pixel_index == 1367) oled_data = 16'b1010110100101001;
    else if (pixel_index == 1368) oled_data = 16'b1010010100101000;
    else if (pixel_index == 1369) oled_data = 16'b1001010010100110;
    else if (pixel_index == 1372 || pixel_index == 2281 || pixel_index == 2376) oled_data = 16'b0101001111000110;
    else if (pixel_index == 1373) oled_data = 16'b0100101111001000;
    else if (pixel_index == 1374 || pixel_index == 1389 || pixel_index == 2477) oled_data = 16'b0101001110000110;
    else if (pixel_index == 1375 || pixel_index == 2773 || pixel_index == 2905) oled_data = 16'b0110001110000011;
    else if (pixel_index == 1376) oled_data = 16'b0110101110000101;
    else if (pixel_index == 1379 || pixel_index == 1461 || pixel_index == 2515) oled_data = 16'b1000010001000111;
    else if (pixel_index == 1381 || pixel_index == 3707) oled_data = 16'b0111001111001110;
    else if (pixel_index == 1382 || pixel_index == 5962) oled_data = 16'b0111110000010000;
    else if (pixel_index == 1383 || pixel_index == 2022 || pixel_index == 2126 || pixel_index == 3026) oled_data = 16'b0110110010110010;
    else if (pixel_index == 1384 || pixel_index == 2217) oled_data = 16'b0101110001010010;
    else if (pixel_index == 1385 || pixel_index == 2265 || pixel_index == 6051) oled_data = 16'b0101101110001111;
    else if (pixel_index == 1392) oled_data = 16'b0011101110000011;
    else if (pixel_index == 1393) oled_data = 16'b0101010000000100;
    else if (pixel_index == 1394) oled_data = 16'b1010111000101110;
    else if (pixel_index == 1395) oled_data = 16'b0110110100100100;
    else if (pixel_index == 1396) oled_data = 16'b1000110110100111;
    else if (pixel_index == 1397) oled_data = 16'b0111101110000110;
    else if (pixel_index == 1398) oled_data = 16'b0010100111000011;
    else if (pixel_index == 1399) oled_data = 16'b0010000111000100;
    else if (pixel_index == 1402) oled_data = 16'b1011010111101100;
    else if (pixel_index == 1403) oled_data = 16'b1010010111100111;
    else if (pixel_index == 1404) oled_data = 16'b1011011001101000;
    else if (pixel_index == 1405) oled_data = 16'b1010010110101101;
    else if (pixel_index == 1406 || pixel_index == 2252) oled_data = 16'b1001110010101011;
    else if (pixel_index == 1408 || pixel_index == 2367 || pixel_index == 2989) oled_data = 16'b0111110001001010;
    else if (pixel_index == 1410 || pixel_index == 2382 || pixel_index == 2904 || pixel_index == 3061) oled_data = 16'b0110001111000101;
    else if (pixel_index == 1411 || pixel_index == 1952) oled_data = 16'b0111110001000111;
    else if (pixel_index == 1413) oled_data = 16'b0111010001000110;
    else if (pixel_index == 1415) oled_data = 16'b1001010101101011;
    else if (pixel_index == 1416 || pixel_index == 2034) oled_data = 16'b0111010011101101;
    else if (pixel_index == 1417 || pixel_index == 2567) oled_data = 16'b0101010001001101;
    else if (pixel_index == 1418 || pixel_index == 2437) oled_data = 16'b0110110010101011;
    else if (pixel_index == 1419 || pixel_index == 2288) oled_data = 16'b0101110000000111;
    else if (pixel_index == 1420) oled_data = 16'b0100101111000111;
    else if (pixel_index == 1423) oled_data = 16'b0111010100100111;
    else if (pixel_index == 1424) oled_data = 16'b0110110010101010;
    else if (pixel_index == 1425 || pixel_index == 2844) oled_data = 16'b0100101111001111;
    else if (pixel_index == 1427) oled_data = 16'b0010101110010100;
    else if (pixel_index == 1428) oled_data = 16'b0011001110010111;
    else if (((pixel_index >= 1429) && (pixel_index <= 1430)) || pixel_index == 1525 || pixel_index == 1620 || pixel_index == 1723 || (pixel_index >= 1725) && (pixel_index <= 1727)) oled_data = 16'b0010001111011001;
    else if (pixel_index == 1431 || pixel_index == 1526 || pixel_index == 1531 || ((pixel_index >= 1629) && (pixel_index <= 1630)) || pixel_index == 1704 || pixel_index == 1711) oled_data = 16'b0001101111011001;
    else if (pixel_index == 1432 || pixel_index == 1440 || pixel_index == 1527 || pixel_index == 1625 || pixel_index == 1710) oled_data = 16'b0001010000011001;
    else if (pixel_index == 1433) oled_data = 16'b0000101111011001;
    else if (pixel_index == 1442) oled_data = 16'b0000101111011000;
    else if (pixel_index == 1443) oled_data = 16'b0000001110011011;
    else if (pixel_index == 1446) oled_data = 16'b0011010000010111;
    else if (pixel_index == 1447 || pixel_index == 1635 || pixel_index == 1920 || pixel_index == 4002) oled_data = 16'b0100110001011000;
    else if (pixel_index == 1448) oled_data = 16'b0101010000010110;
    else if (pixel_index == 1449) oled_data = 16'b0111010011110000;
    else if (pixel_index == 1450 || pixel_index == 2046 || pixel_index == 2442 || pixel_index == 2722) oled_data = 16'b1000110011101101;
    else if (pixel_index == 1451 || pixel_index == 3160) oled_data = 16'b1001010011101001;
    else if (pixel_index == 1452) oled_data = 16'b1010110101101010;
    else if (pixel_index == 1453) oled_data = 16'b1010110110101000;
    else if (pixel_index == 1454 || pixel_index == 2340) oled_data = 16'b1010010101100101;
    else if (pixel_index == 1457) oled_data = 16'b1000110011100110;
    else if (((pixel_index >= 1458) && (pixel_index <= 1459)) || pixel_index == 1470 || pixel_index == 2615) oled_data = 16'b1000110011100101;
    else if (pixel_index == 1460 || pixel_index == 1865) oled_data = 16'b1000010010100101;
    else if (pixel_index == 1462 || pixel_index == 1782) oled_data = 16'b1000110011101000;
    else if (pixel_index == 1463) oled_data = 16'b1000010011101000;
    else if (pixel_index == 1464 || pixel_index == 1597 || pixel_index == 2768) oled_data = 16'b0111010010100111;
    else if (pixel_index == 1465 || ((pixel_index >= 1558) && (pixel_index <= 1559)) || pixel_index == 2286 || pixel_index == 2775 || pixel_index == 2958) oled_data = 16'b0111010000000110;
    else if (pixel_index == 1466 || pixel_index == 1857 || pixel_index == 2057) oled_data = 16'b1000010000000110;
    else if (pixel_index == 1467 || pixel_index == 2050) oled_data = 16'b1000110010100100;
    else if (pixel_index == 1468) oled_data = 16'b1001110100100110;
    else if (pixel_index == 1472) oled_data = 16'b0111110001000110;
    else if (pixel_index == 1473 || pixel_index == 1997 || pixel_index == 2996) oled_data = 16'b0111010001000100;
    else if (pixel_index == 1474 || pixel_index == 1546 || pixel_index == 1564) oled_data = 16'b1001010010101000;
    else if (pixel_index == 1477 || pixel_index == 1979 || pixel_index == 2895) oled_data = 16'b0110010000000111;
    else if (pixel_index == 1481 || pixel_index == 3654) oled_data = 16'b0111010001001100;
    else if (pixel_index == 1482 || pixel_index == 3229) oled_data = 16'b0101101101001001;
    else if (pixel_index == 1483) oled_data = 16'b0101101100001010;
    else if (pixel_index == 1484 || pixel_index == 2639) oled_data = 16'b0110001101001001;
    else if (pixel_index == 1487 || pixel_index == 2082) oled_data = 16'b0011001010000010;
    else if (pixel_index == 1488) oled_data = 16'b0001100101000010;
    else if (pixel_index == 1490 || pixel_index == 2907) oled_data = 16'b1000110010101011;
    else if (pixel_index == 1496) oled_data = 16'b1001110111101010;
    else if (pixel_index == 1497) oled_data = 16'b1010111000101010;
    else if (pixel_index == 1498) oled_data = 16'b1101011010101101;
    else if (pixel_index == 1501 || pixel_index == 3161) oled_data = 16'b1001110101101100;
    else if (pixel_index == 1502) oled_data = 16'b1010110110101010;
    else if (pixel_index == 1503 || pixel_index == 1506 || pixel_index == 2808) oled_data = 16'b0110010000000100;
    else if (pixel_index == 1504 || pixel_index == 1553 || pixel_index == 1590 || pixel_index == 2672) oled_data = 16'b0110110001000111;
    else if (pixel_index == 1505 || pixel_index == 1884) oled_data = 16'b0101101111000101;
    else if (pixel_index == 1510 || pixel_index == 1783) oled_data = 16'b1000010100101010;
    else if (pixel_index == 1511 || pixel_index == 2150) oled_data = 16'b1000110100101101;
    else if (pixel_index == 1512 || pixel_index == 1542 || pixel_index == 2195 || pixel_index == 3992) oled_data = 16'b0101110001010001;
    else if (pixel_index == 1513) oled_data = 16'b0011110000010010;
    else if (pixel_index == 1514 || pixel_index == 1521) oled_data = 16'b0100010000010010;
    else if (pixel_index == 1515 || pixel_index == 1790) oled_data = 16'b0100010000001111;
    else if (pixel_index == 1516) oled_data = 16'b0100101111001101;
    else if (pixel_index == 1517) oled_data = 16'b0100101111001110;
    else if (pixel_index == 1518 || pixel_index == 2027) oled_data = 16'b0100110000001111;
    else if (pixel_index == 1520 || pixel_index == 3222) oled_data = 16'b0110110001010001;
    else if (pixel_index == 1522) oled_data = 16'b0011101110010010;
    else if (pixel_index == 1523) oled_data = 16'b0011101110010100;
    else if (pixel_index == 1524 || pixel_index == 1539) oled_data = 16'b0010101111011000;
    else if (pixel_index == 1528) oled_data = 16'b0001110000011000;
    else if (pixel_index == 1529) oled_data = 16'b0010001111011000;
    else if (pixel_index == 1532 || pixel_index == 3920) oled_data = 16'b0001101111011000;
    else if (pixel_index == 1536) oled_data = 16'b0001010001011011;
    else if (pixel_index == 1538 || pixel_index == 1621 || pixel_index == 1626 || pixel_index == 1721) oled_data = 16'b0001101111011010;
    else if (pixel_index == 1540 || ((pixel_index >= 1610) && (pixel_index <= 1611)) || pixel_index == 1617) oled_data = 16'b0010101111010111;
    else if (pixel_index == 1541 || pixel_index == 2223) oled_data = 16'b0100110000010100;
    else if (pixel_index == 1543 || pixel_index == 2866) oled_data = 16'b0110110010101110;
    else if (pixel_index == 1544 || pixel_index == 2968) oled_data = 16'b0111110010101011;
    else if (pixel_index == 1545 || pixel_index == 1847 || pixel_index == 3064) oled_data = 16'b0111110001001001;
    else if (pixel_index == 1549 || pixel_index == 2613) oled_data = 16'b1001010011100110;
    else if (pixel_index == 1550 || pixel_index == 1957 || pixel_index == 2055 || pixel_index == 2423 || pixel_index == 2812) oled_data = 16'b1000010010101000;
    else if (pixel_index == 1551 || pixel_index == 1740 || pixel_index == 1772 || pixel_index == 2420 || pixel_index == 2872) oled_data = 16'b0111010010101011;
    else if (pixel_index == 1552) oled_data = 16'b0110110010101001;
    else if (pixel_index == 1554 || pixel_index == 2375) oled_data = 16'b0110001111000100;
    else if (pixel_index == 1555 || pixel_index == 2087 || pixel_index == 2186) oled_data = 16'b0101101110000011;
    else if (pixel_index == 1556 || pixel_index == 1671 || pixel_index == 1777 || pixel_index == 2862) oled_data = 16'b0110001111000110;
    else if (pixel_index == 1557 || pixel_index == 1892 || pixel_index == 2289 || pixel_index == 2341) oled_data = 16'b0110010001001000;
    else if (pixel_index == 1565) oled_data = 16'b1000010001000011;
    else if (pixel_index == 1566 || pixel_index == 2189) oled_data = 16'b0111110000000011;
    else if (pixel_index == 1569 || pixel_index == 2711) oled_data = 16'b0111110010100100;
    else if (pixel_index == 1571) oled_data = 16'b1010010011100111;
    else if (pixel_index == 1572) oled_data = 16'b1001110010100111;
    else if (pixel_index == 1573 || pixel_index == 1751 || pixel_index == 3062) oled_data = 16'b0110101111000101;
    else if (pixel_index == 1575) oled_data = 16'b0101001111000111;
    else if (pixel_index == 1578 || pixel_index == 2868 || pixel_index == 2964) oled_data = 16'b0101101111001000;
    else if (pixel_index == 1579 || pixel_index == 3558) oled_data = 16'b0110101111001011;
    else if (pixel_index == 1580) oled_data = 16'b0110101110001011;
    else if (pixel_index == 1583 || pixel_index == 1984) oled_data = 16'b0011101011000010;
    else if (pixel_index == 1585) oled_data = 16'b0000100100000001;
    else if (pixel_index == 1586) oled_data = 16'b0001100111000100;
    else if (pixel_index == 1587 || pixel_index == 2730) oled_data = 16'b0011001001000011;
    else if (pixel_index == 1589 || pixel_index == 2823 || pixel_index == 3360) oled_data = 16'b0101101100000110;
    else if (pixel_index == 1591) oled_data = 16'b1001110111101001;
    else if (pixel_index == 1593) oled_data = 16'b1010010111101001;
    else if (pixel_index == 1594) oled_data = 16'b1011111000101101;
    else if (pixel_index == 1595 || pixel_index == 1739 || pixel_index == 2245) oled_data = 16'b1000010100101011;
    else if (pixel_index == 1596) oled_data = 16'b0111110011101011;
    else if (pixel_index == 1598) oled_data = 16'b1001110010101010;
    else if (pixel_index == 1599 || pixel_index == 1691 || pixel_index == 2871) oled_data = 16'b0111010001001001;
    else if (pixel_index == 1600) oled_data = 16'b0110010010101000;
    else if (((pixel_index >= 1601) && (pixel_index <= 1603)) || pixel_index == 1894) oled_data = 16'b0111010011101000;
    else if (pixel_index == 1604 || pixel_index == 1900 || pixel_index == 2999) oled_data = 16'b0111010010101001;
    else if (pixel_index == 1605 || pixel_index == 1836 || pixel_index == 2679) oled_data = 16'b0110010001001100;
    else if (pixel_index == 1606 || pixel_index == 2770 || pixel_index == 2984 || pixel_index == 3993) oled_data = 16'b0110010000001110;
    else if (pixel_index == 1608 || pixel_index == 1728) oled_data = 16'b0100010001010100;
    else if (pixel_index == 1609 || pixel_index == 1794 || pixel_index == 2592) oled_data = 16'b0011010000010110;
    else if (pixel_index == 1612) oled_data = 16'b0011010000010101;
    else if (pixel_index == 1613) oled_data = 16'b0100110001010100;
    else if (pixel_index == 1614) oled_data = 16'b0100110000010110;
    else if (pixel_index == 1615 || pixel_index == 4004) oled_data = 16'b0011110000010111;
    else if (pixel_index == 1616) oled_data = 16'b0100001111010111;
    else if (pixel_index == 1618 || pixel_index == 2400) oled_data = 16'b0010101111010110;
    else if (((pixel_index >= 1623) && (pixel_index <= 1624)) || pixel_index == 1722) oled_data = 16'b0001110000011001;
    else if (pixel_index == 1631) oled_data = 16'b0010001110011001;
    else if (pixel_index == 1632 || pixel_index == 1701) oled_data = 16'b0100010000010011;
    else if (pixel_index == 1634) oled_data = 16'b0100110000010111;
    else if (pixel_index == 1636 || (pixel_index >= 4000) && (pixel_index <= 4001)) oled_data = 16'b0101010010111000;
    else if (pixel_index == 1637 || pixel_index == 4705) oled_data = 16'b0111110010110011;
    else if (pixel_index == 1639) oled_data = 16'b1001110011100111;
    else if (pixel_index == 1640) oled_data = 16'b1001110011100101;
    else if (pixel_index == 1641 || pixel_index == 1690) oled_data = 16'b1001010010100111;
    else if (pixel_index == 1645 || pixel_index == 2000 || pixel_index == 2053 || pixel_index == 2706) oled_data = 16'b1000110011101001;
    else if (pixel_index == 1646 || pixel_index == 2267 || pixel_index == 2365) oled_data = 16'b0111110010101010;
    else if (pixel_index == 1650) oled_data = 16'b0100101111000101;
    else if (pixel_index == 1652 || pixel_index == 1787) oled_data = 16'b0101101111000111;
    else if (pixel_index == 1656 || pixel_index == 1688 || pixel_index == 2095 || pixel_index == 2671 || (pixel_index >= 2809) && (pixel_index <= 2810)) oled_data = 16'b0110110000000100;
    else if (pixel_index == 1657 || pixel_index == 2427 || pixel_index == 2708) oled_data = 16'b1000010011100110;
    else if (pixel_index == 1660 || pixel_index == 1754) oled_data = 16'b1000010001001000;
    else if (((pixel_index >= 1661) && (pixel_index <= 1662)) || pixel_index == 1763) oled_data = 16'b1000010000000100;
    else if (pixel_index == 1663) oled_data = 16'b0111110000000010;
    else if (pixel_index == 1664 || pixel_index == 2619) oled_data = 16'b0111110001000011;
    else if (pixel_index == 1665) oled_data = 16'b1000010010100011;
    else if (pixel_index == 1666 || pixel_index == 1954) oled_data = 16'b1000010001000010;
    else if (pixel_index == 1667) oled_data = 16'b1001110001000101;
    else if (pixel_index == 1668) oled_data = 16'b1001110010100110;
    else if (pixel_index == 1669 || pixel_index == 1768 || pixel_index == 2075 || pixel_index == 2906) oled_data = 16'b0111001111000100;
    else if (pixel_index == 1670 || pixel_index == 2863) oled_data = 16'b0111010000000101;
    else if (pixel_index == 1673 || pixel_index == 2967) oled_data = 16'b0111010000001001;
    else if (pixel_index == 1674 || pixel_index == 3001) oled_data = 16'b0110101111001000;
    else if (pixel_index == 1676 || pixel_index == 1835 || pixel_index == 2771 || pixel_index == 2916) oled_data = 16'b0110010001001011;
    else if (pixel_index == 1677) oled_data = 16'b0100101111001011;
    else if (pixel_index == 1678) oled_data = 16'b0101101110001001;
    else if (pixel_index == 1679) oled_data = 16'b0100001101000100;
    else if (pixel_index == 1681) oled_data = 16'b0010100111000001;
    else if (pixel_index == 1682) oled_data = 16'b0000100101000010;
    else if (pixel_index == 1683) oled_data = 16'b0001100111000000;
    else if (pixel_index == 1686) oled_data = 16'b0111110100100111;
    else if (pixel_index == 1687) oled_data = 16'b1001010111101000;
    else if (pixel_index == 1689) oled_data = 16'b1000110010101010;
    else if (pixel_index == 1692 || pixel_index == 1901 || pixel_index == 2669) oled_data = 16'b0110110001001001;
    else if (pixel_index == 1695 || pixel_index == 2764) oled_data = 16'b0110010010101100;
    else if (pixel_index == 1696) oled_data = 16'b0101110001001011;
    else if (pixel_index == 1697 || pixel_index == 1942 || pixel_index == 2025 || pixel_index == 2867) oled_data = 16'b0110010010101110;
    else if (((pixel_index >= 1698) && (pixel_index <= 1699)) || pixel_index == 1887 || pixel_index == 2569) oled_data = 16'b0101010001001111;
    else if (pixel_index == 1700) oled_data = 16'b0100110001010000;
    else if (pixel_index == 1703) oled_data = 16'b0010110000010111;
    else if (pixel_index == 1707) oled_data = 16'b0000110000011011;
    else if (pixel_index == 1708 || pixel_index == 1717 || pixel_index == 1806 || pixel_index == 1813) oled_data = 16'b0001010000011010;
    else if (pixel_index == 1709 || pixel_index == 1807 || pixel_index == 1822) oled_data = 16'b0010010000011001;
    else if (pixel_index == 1712) oled_data = 16'b0001101110011010;
    else if (pixel_index == 1713 || pixel_index == 1809 || pixel_index == 1812) oled_data = 16'b0001010000011011;
    else if (pixel_index == 1714) oled_data = 16'b0001001111011010;
    else if (pixel_index == 1715) oled_data = 16'b0001001110011010;
    else if (pixel_index == 1716) oled_data = 16'b0001001111011011;
    else if (pixel_index == 1718 || pixel_index == 1814 || pixel_index == 1816 || pixel_index == 1818 || pixel_index == 1820 || pixel_index == 1823) oled_data = 16'b0010010000011010;
    else if (pixel_index == 1724 || pixel_index == 1821) oled_data = 16'b0010001111011010;
    else if (pixel_index == 1730) oled_data = 16'b0101110000010100;
    else if (pixel_index == 1731 || pixel_index == 4707 || pixel_index == 6008 || pixel_index == 6103) oled_data = 16'b1000010001010010;
    else if (pixel_index == 1732 || pixel_index == 2249 || pixel_index == 3080) oled_data = 16'b1000010001010000;
    else if (pixel_index == 1733) oled_data = 16'b1001110011101111;
    else if (pixel_index == 1734 || pixel_index == 3179) oled_data = 16'b1010010100101100;
    else if (pixel_index == 1735) oled_data = 16'b1010110101101001;
    else if (pixel_index == 1738) oled_data = 16'b1000010011101011;
    else if (pixel_index == 1744 || pixel_index == 1784 || pixel_index == 2965) oled_data = 16'b0101101110000101;
    else if (pixel_index == 1746 || pixel_index == 1937) oled_data = 16'b0011101011000100;
    else if (pixel_index == 1747 || pixel_index == 3225 || pixel_index == 3936) oled_data = 16'b0100001100000111;
    else if (pixel_index == 1748 || pixel_index == 1883) oled_data = 16'b0101010000001001;
    else if (pixel_index == 1749 || pixel_index == 2769 || pixel_index == 2894) oled_data = 16'b0101110000001011;
    else if (pixel_index == 1752 || pixel_index == 1770) oled_data = 16'b0111110010101000;
    else if (pixel_index == 1756) oled_data = 16'b0111110000000111;
    else if (pixel_index == 1758) oled_data = 16'b1001010001000011;
    else if (pixel_index == 1759) oled_data = 16'b1000010010100010;
    else if (pixel_index == 1760) oled_data = 16'b1000110010100001;
    else if (pixel_index == 1761 || pixel_index == 1959 || pixel_index == 1999 || pixel_index == 2713 || pixel_index == 2716 || pixel_index == 2899) oled_data = 16'b1000110010100101;
    else if (pixel_index == 1764 || pixel_index == 1861 || pixel_index == 2047) oled_data = 16'b1000110000000101;
    else if (pixel_index == 1765) oled_data = 16'b1000001110000010;
    else if (pixel_index == 1766) oled_data = 16'b0111001110000010;
    else if (pixel_index == 1767) oled_data = 16'b0111101110000011;
    else if (pixel_index == 1769 || pixel_index == 2348) oled_data = 16'b1000110010101000;
    else if (pixel_index == 1771) oled_data = 16'b1001010100101010;
    else if (pixel_index == 1774) oled_data = 16'b0110101110001010;
    else if (pixel_index == 1775 || pixel_index == 1969) oled_data = 16'b0110001100000110;
    else if (pixel_index == 1776 || pixel_index == 2032 || pixel_index == 2966) oled_data = 16'b0110001110000110;
    else if (pixel_index == 1778) oled_data = 16'b0010000110000001;
    else if (pixel_index == 1779) oled_data = 16'b0010001000000010;
    else if (pixel_index == 1780 || pixel_index == 2268 || pixel_index == 2371) oled_data = 16'b0111010001001000;
    else if (pixel_index == 1781 || pixel_index == 1877) oled_data = 16'b1011011001101100;
    else if (pixel_index == 1785 || pixel_index == 2820) oled_data = 16'b0110001101000100;
    else if (pixel_index == 1788) oled_data = 16'b0110010001000111;
    else if (pixel_index == 1789 || pixel_index == 2377) oled_data = 16'b0101110000001001;
    else if (pixel_index == 1791) oled_data = 16'b0101010010110001;
    else if (pixel_index == 1792) oled_data = 16'b0011110000010011;
    else if (pixel_index == 1793 || pixel_index == 3896) oled_data = 16'b0011110001010101;
    else if (pixel_index == 1796 || pixel_index == 2123 || pixel_index == 2888) oled_data = 16'b0100010010110101;
    else if (pixel_index == 1797 || pixel_index == 2133) oled_data = 16'b0100010010110110;
    else if (pixel_index == 1798 || pixel_index == 2305) oled_data = 16'b0011010001010110;
    else if (pixel_index == 1799 || pixel_index == 2306 || pixel_index == 2326) oled_data = 16'b0011010010110111;
    else if (pixel_index == 1800) oled_data = 16'b0011010010111000;
    else if (pixel_index == 1801 || pixel_index == 2100 || pixel_index == 2137) oled_data = 16'b0011110010111000;
    else if (((pixel_index >= 1802) && (pixel_index <= 1803)) || pixel_index == 4009) oled_data = 16'b0010010001011000;
    else if (pixel_index == 1804) oled_data = 16'b0001010001011001;
    else if (pixel_index == 1808 || pixel_index == 1914 || pixel_index == 1917) oled_data = 16'b0001110001011011;
    else if ((pixel_index >= 1810) && (pixel_index <= 1811)) oled_data = 16'b0001010000011100;
    else if (pixel_index == 1824) oled_data = 16'b0011010000011001;
    else if (pixel_index == 1825) oled_data = 16'b0100010000011000;
    else if (pixel_index == 1826) oled_data = 16'b0110010010110011;
    else if (pixel_index == 1827 || pixel_index == 1923 || pixel_index == 3655) oled_data = 16'b1000010001001100;
    else if (pixel_index == 1828) oled_data = 16'b1001010000001011;
    else if (pixel_index == 1829) oled_data = 16'b1010010011101101;
    else if (pixel_index == 1830 || pixel_index == 2145) oled_data = 16'b1001010100110000;
    else if (pixel_index == 1831) oled_data = 16'b1001110101101110;
    else if (pixel_index == 1833) oled_data = 16'b0111010100110000;
    else if (pixel_index == 1838) oled_data = 16'b0101110010101111;
    else if (pixel_index == 1839) oled_data = 16'b0101001110001001;
    else if (pixel_index == 1841 || pixel_index == 3227 || pixel_index == 3554) oled_data = 16'b0011101001000001;
    else if (pixel_index == 1843 || pixel_index == 2481) oled_data = 16'b0101001111001011;
    else if (pixel_index == 1844 || pixel_index == 2979) oled_data = 16'b0101110001001100;
    else if (pixel_index == 1845) oled_data = 16'b0101110000001010;
    else if (pixel_index == 1849 || pixel_index == 2721) oled_data = 16'b1000010010101010;
    else if (((pixel_index >= 1850) && (pixel_index <= 1851)) || pixel_index == 2801 || pixel_index == 3054) oled_data = 16'b1000010001001001;
    else if (pixel_index == 1852 || pixel_index == 3002 || pixel_index == 3153) oled_data = 16'b0111101111001000;
    else if (pixel_index == 1854) oled_data = 16'b1001010010100101;
    else if (pixel_index == 1855) oled_data = 16'b1000110001000011;
    else if (pixel_index == 1856) oled_data = 16'b1000110001000101;
    else if (pixel_index == 1858 || pixel_index == 1992) oled_data = 16'b0101101111000011;
    else if (pixel_index == 1862) oled_data = 16'b0111101111000010;
    else if (pixel_index == 1863) oled_data = 16'b0111101111000001;
    else if (pixel_index == 1864) oled_data = 16'b1000110010100010;
    else if (pixel_index == 1866) oled_data = 16'b0111101111000100;
    else if (((pixel_index >= 1869) && (pixel_index <= 1870)) || pixel_index == 3057) oled_data = 16'b0110001111001011;
    else if (pixel_index == 1871 || pixel_index == 2724) oled_data = 16'b0111001111001010;
    else if (pixel_index == 1872) oled_data = 16'b0111101111001010;
    else if (pixel_index == 1873) oled_data = 16'b1000010000001001;
    else if (pixel_index == 1874) oled_data = 16'b0100000110000010;
    else if (pixel_index == 1875 || pixel_index == 2081 || pixel_index == 3323) oled_data = 16'b0011101010000010;
    else if (pixel_index == 1879 || pixel_index == 3321) oled_data = 16'b0101101101001010;
    else if (pixel_index == 1881 || pixel_index == 2085) oled_data = 16'b0100101100000001;
    else if (pixel_index == 1882) oled_data = 16'b0100110000000101;
    else if (pixel_index == 1886 || pixel_index == 4129) oled_data = 16'b0101010000001011;
    else if (pixel_index == 1888) oled_data = 16'b0011001110001100;
    else if (pixel_index == 1889) oled_data = 16'b0011001110001011;
    else if (pixel_index == 1890) oled_data = 16'b0100101110001011;
    else if (pixel_index == 1893 || pixel_index == 2096) oled_data = 16'b0111010010101000;
    else if (pixel_index == 1895 || pixel_index == 1897) oled_data = 16'b1000110100101000;
    else if (pixel_index == 1899 || pixel_index == 2525) oled_data = 16'b0111110011101000;
    else if (pixel_index == 1902 || pixel_index == 2725) oled_data = 16'b0110110000001010;
    else if (pixel_index == 1903 || pixel_index == 2961) oled_data = 16'b0111010011101100;
    else if (pixel_index == 1904) oled_data = 16'b0110010011110000;
    else if (pixel_index == 1905 || pixel_index == 3748) oled_data = 16'b0101010011110010;
    else if (pixel_index == 1906) oled_data = 16'b0100110010110100;
    else if (pixel_index == 1907 || pixel_index == 2131 || pixel_index == 2221) oled_data = 16'b0011110010110111;
    else if (pixel_index == 1908 || pixel_index == 2006) oled_data = 16'b0010110001011001;
    else if (pixel_index == 1909 || pixel_index == 2007) oled_data = 16'b0010110001011010;
    else if (pixel_index == 1910) oled_data = 16'b0001110010111011;
    else if (pixel_index == 1911) oled_data = 16'b0001110010111010;
    else if (pixel_index == 1912) oled_data = 16'b0001110001011010;
    else if (pixel_index == 1913) oled_data = 16'b0010010001011010;
    else if (pixel_index == 1915) oled_data = 16'b0001110000011011;
    else if (pixel_index == 1918 || ((pixel_index >= 2010) && (pixel_index <= 2011)) || (pixel_index >= 2014) && (pixel_index <= 2015)) oled_data = 16'b0010010001011011;
    else if (pixel_index == 1919) oled_data = 16'b0010010000011011;
    else if (pixel_index == 1921 || pixel_index == 2138) oled_data = 16'b0101010010110111;
    else if (pixel_index == 1924 || pixel_index == 2421 || pixel_index == 2800 || pixel_index == 3519) oled_data = 16'b0111110001001011;
    else if (pixel_index == 1925) oled_data = 16'b1000010010101111;
    else if ((pixel_index >= 1927) && (pixel_index <= 1928)) oled_data = 16'b0111010011110011;
    else if (pixel_index == 1929 || pixel_index == 2019 || pixel_index == 2218 || pixel_index == 2858 || pixel_index == 3106) oled_data = 16'b0110110010110001;
    else if (pixel_index == 1930) oled_data = 16'b0110110000001101;
    else if (pixel_index == 1931 || pixel_index == 2253 || pixel_index == 2290) oled_data = 16'b0110110000001011;
    else if (pixel_index == 1933 || pixel_index == 2473) oled_data = 16'b0101110001001101;
    else if (pixel_index == 1934 || pixel_index == 2665) oled_data = 16'b0101010010110000;
    else if (pixel_index == 1935) oled_data = 16'b0100101101000111;
    else if (pixel_index == 1939) oled_data = 16'b0111010010101111;
    else if (pixel_index == 1941 || pixel_index == 2463 || pixel_index == 2963) oled_data = 16'b0111010010101101;
    else if (pixel_index == 1943 || pixel_index == 2122 || pixel_index == 2342) oled_data = 16'b0110010010110000;
    else if (pixel_index == 1945 || pixel_index == 2817) oled_data = 16'b1000010010101110;
    else if (pixel_index == 1946) oled_data = 16'b0111110001001101;
    else if (pixel_index == 1948 || pixel_index == 1972 || pixel_index == 2512 || pixel_index == 3189) oled_data = 16'b1001010010101010;
    else if (pixel_index == 1951) oled_data = 16'b1000010000000101;
    else if (pixel_index == 1953) oled_data = 16'b0110110001000100;
    else if (pixel_index == 1955 || pixel_index == 2611) oled_data = 16'b0111110000000101;
    else if (pixel_index == 1956) oled_data = 16'b1001010001001000;
    else if (pixel_index == 1960) oled_data = 16'b1001110010100010;
    else if (pixel_index == 1961) oled_data = 16'b1000110000000011;
    else if (pixel_index == 1962) oled_data = 16'b0111101101000010;
    else if (pixel_index == 1963) oled_data = 16'b0111101110000010;
    else if (pixel_index == 1964) oled_data = 16'b0110101101000110;
    else if (pixel_index == 1965 || pixel_index == 2564) oled_data = 16'b0101101111001110;
    else if (pixel_index == 1966) oled_data = 16'b0101001111010001;
    else if (pixel_index == 1967) oled_data = 16'b1001010010110001;
    else if (pixel_index == 1968 || pixel_index == 2255) oled_data = 16'b1000101110001010;
    else if (pixel_index == 1970) oled_data = 16'b0111001101000110;
    else if (pixel_index == 1971) oled_data = 16'b1000001100001000;
    else if (pixel_index == 1973 || pixel_index == 3255) oled_data = 16'b1001110101101101;
    else if (pixel_index == 1974 || pixel_index == 2824) oled_data = 16'b0101001111001101;
    else if (pixel_index == 1975) oled_data = 16'b0011101100001101;
    else if (pixel_index == 1980 || pixel_index == 2573 || pixel_index == 2869) oled_data = 16'b0101101110000111;
    else if (pixel_index == 1981) oled_data = 16'b0110101101000101;
    else if (pixel_index == 1983 || pixel_index == 3228) oled_data = 16'b0100001010000100;
    else if (pixel_index == 1986) oled_data = 16'b0100101010000010;
    else if (pixel_index == 1987) oled_data = 16'b0110001101000010;
    else if (pixel_index == 1988) oled_data = 16'b0101101101000001;
    else if (pixel_index == 1989) oled_data = 16'b0100101110000010;
    else if (pixel_index == 1990) oled_data = 16'b0100101111000010;
    else if (pixel_index == 1991 || pixel_index == 2901) oled_data = 16'b0110001111000010;
    else if (pixel_index == 1993) oled_data = 16'b0110110001000011;
    else if (pixel_index == 1995 || pixel_index == 2089) oled_data = 16'b0110010000000011;
    else if (pixel_index == 1996) oled_data = 16'b0110110000000011;
    else if (pixel_index == 1998 || pixel_index == 2767) oled_data = 16'b1000010001000100;
    else if (pixel_index == 2001 || pixel_index == 2097) oled_data = 16'b0111010011101010;
    else if (pixel_index == 2002) oled_data = 16'b0111010011101110;
    else if (pixel_index == 2003 || pixel_index == 2043 || pixel_index == 2247) oled_data = 16'b0111110011110000;
    else if (pixel_index == 2004 || pixel_index == 2919) oled_data = 16'b0110010011110101;
    else if (pixel_index == 2005 || pixel_index == 2136 || pixel_index == 2389) oled_data = 16'b0100010010111000;
    else if (pixel_index == 2008) oled_data = 16'b0010110010111010;
    else if (pixel_index == 2009 || pixel_index == 2102 || ((pixel_index >= 2104) && (pixel_index <= 2105)) || ((pixel_index >= 2108) && (pixel_index <= 2110)) || pixel_index == 2198 || pixel_index == 2235 || pixel_index == 2295) oled_data = 16'b0010110010111011;
    else if (((pixel_index >= 2012) && (pixel_index <= 2013)) || pixel_index == 2107 || pixel_index == 2202 || pixel_index == 2232) oled_data = 16'b0010010010111011;
    else if (pixel_index == 2016 || pixel_index == 3119 || pixel_index == 4996) oled_data = 16'b0110001110010000;
    else if (pixel_index == 2017 || pixel_index == 2114) oled_data = 16'b0110110000010001;
    else if (pixel_index == 2018) oled_data = 16'b0111110010110010;
    else if (pixel_index == 2021 || pixel_index == 3365 || pixel_index == 3505) oled_data = 16'b0111010010110011;
    else if (pixel_index == 2023) oled_data = 16'b0110010001010010;
    else if (pixel_index == 2029 || pixel_index == 2388) oled_data = 16'b0101110010110010;
    else if (pixel_index == 2030 || pixel_index == 2980) oled_data = 16'b0101110010110001;
    else if (pixel_index == 2031) oled_data = 16'b0101101110001000;
    else if (pixel_index == 2035 || pixel_index == 3319) oled_data = 16'b0111010100110011;
    else if ((pixel_index >= 2038) && (pixel_index <= 2039)) oled_data = 16'b0110010100110100;
    else if (pixel_index == 2040) oled_data = 16'b0110010011110100;
    else if (pixel_index == 2042 || pixel_index == 2418 || pixel_index == 2723 || pixel_index == 3651) oled_data = 16'b0111010010110001;
    else if (pixel_index == 2044 || pixel_index == 3560) oled_data = 16'b0111110010110000;
    else if (pixel_index == 2045) oled_data = 16'b1000010100110001;
    else if (pixel_index == 2048) oled_data = 16'b1000110001001000;
    else if (pixel_index == 2049 || pixel_index == 2424) oled_data = 16'b1000110010100111;
    else if (pixel_index == 2056 || pixel_index == 2705) oled_data = 16'b1000110001000111;
    else if (pixel_index == 2058) oled_data = 16'b0111001100000101;
    else if (pixel_index == 2059) oled_data = 16'b0111001100000011;
    else if (pixel_index == 2060 || pixel_index == 2870) oled_data = 16'b0110101110000110;
    else if (pixel_index == 2061) oled_data = 16'b0101001111010010;
    else if (pixel_index == 2064) oled_data = 16'b0111001101001100;
    else if (pixel_index == 2065) oled_data = 16'b0110001001001000;
    else if (pixel_index == 2066) oled_data = 16'b0101101001001001;
    else if (pixel_index == 2067 || pixel_index == 3024) oled_data = 16'b0100100111000110;
    else if (pixel_index == 2068) oled_data = 16'b0101101010001001;
    else if (pixel_index == 2070 || pixel_index == 2165) oled_data = 16'b0101001101001110;
    else if (pixel_index == 2071) oled_data = 16'b0100101010001010;
    else if (pixel_index == 2073) oled_data = 16'b0101101101000111;
    else if (pixel_index == 2074) oled_data = 16'b1000001110000100;
    else if (pixel_index == 2076) oled_data = 16'b0101001100000001;
    else if (pixel_index == 2077 || pixel_index == 2086 || pixel_index == 2172) oled_data = 16'b0101001101000010;
    else if (pixel_index == 2078) oled_data = 16'b0101001111000100;
    else if (pixel_index == 2083 || pixel_index == 3419) oled_data = 16'b0100001100000011;
    else if (pixel_index == 2084) oled_data = 16'b0100101100000011;
    else if (pixel_index == 2090 || (pixel_index >= 2187) && (pixel_index <= 2188)) oled_data = 16'b0110101111000011;
    else if (pixel_index == 2091 || pixel_index == 2370) oled_data = 16'b0110101111000100;
    else if (pixel_index == 2098) oled_data = 16'b0110110010101111;
    else if (pixel_index == 2099 || pixel_index == 3806) oled_data = 16'b0101010010110011;
    else if (pixel_index == 2101) oled_data = 16'b0011010001011011;
    else if (pixel_index == 2103 || pixel_index == 2229 || pixel_index == 2318 || pixel_index == 2406) oled_data = 16'b0010010010111100;
    else if (pixel_index == 2106 || pixel_index == 2225 || (pixel_index >= 2407) && (pixel_index <= 2408)) oled_data = 16'b0010110010111100;
    else if (pixel_index == 2111 || pixel_index == 2203) oled_data = 16'b0010110001011011;
    else if (pixel_index == 2113) oled_data = 16'b0110001101001010;
    else if (pixel_index == 2116 || pixel_index == 4418) oled_data = 16'b0111010011110110;
    else if (pixel_index == 2117) oled_data = 16'b0111010011110100;
    else if (pixel_index == 2118) oled_data = 16'b0110010001010000;
    else if (pixel_index == 2119 || pixel_index == 3997) oled_data = 16'b0101110000010001;
    else if (pixel_index == 2124) oled_data = 16'b0110010100110010;
    else if (pixel_index == 2125 || pixel_index == 2788) oled_data = 16'b0100110011110110;
    else if (pixel_index == 2127 || pixel_index == 3223) oled_data = 16'b0110001111001101;
    else if (pixel_index == 2128) oled_data = 16'b0110101111001101;
    else if (pixel_index == 2130) oled_data = 16'b0101010011110101;
    else if (pixel_index == 2132 || pixel_index == 3169) oled_data = 16'b0110010010110110;
    else if (pixel_index == 2134) oled_data = 16'b0011110011111001;
    else if (pixel_index == 2135 || pixel_index == 2416 || pixel_index == 2787) oled_data = 16'b0100110011111001;
    else if (pixel_index == 2139 || pixel_index == 2315) oled_data = 16'b0100110010110111;
    else if (pixel_index == 2140) oled_data = 16'b0100010001010111;
    else if (pixel_index == 2141 || pixel_index == 3809) oled_data = 16'b0101010010111001;
    else if (pixel_index == 2142 || pixel_index == 4417) oled_data = 16'b0111010010110101;
    else if (pixel_index == 2143 || pixel_index == 2156) oled_data = 16'b0111110000001010;
    else if (pixel_index == 2146 || pixel_index == 3559) oled_data = 16'b0111110010101110;
    else if (pixel_index == 2147 || pixel_index == 3003) oled_data = 16'b1000010011101111;
    else if (pixel_index == 2148) oled_data = 16'b1000010101101110;
    else if (pixel_index == 2149) oled_data = 16'b1001010100101101;
    else if (pixel_index == 2152) oled_data = 16'b1000001111001100;
    else if (pixel_index == 2154) oled_data = 16'b0110001100001011;
    else if (pixel_index == 2155 || pixel_index == 2930) oled_data = 16'b0110101101001001;
    else if (pixel_index == 2157) oled_data = 16'b0011010000010011;
    else if (pixel_index == 2160) oled_data = 16'b1001010000001111;
    else if (pixel_index == 2161) oled_data = 16'b1001110001010000;
    else if (pixel_index == 2162) oled_data = 16'b0111001011001110;
    else if (pixel_index == 2163) oled_data = 16'b0010000100000011;
    else if (pixel_index == 2164) oled_data = 16'b0011000110000110;
    else if (pixel_index == 2166) oled_data = 16'b0101101101001101;
    else if (pixel_index == 2167) oled_data = 16'b0110001011001000;
    else if (pixel_index == 2168) oled_data = 16'b0110101011001010;
    else if (pixel_index == 2169) oled_data = 16'b0110001110001011;
    else if (pixel_index == 2170 || pixel_index == 2959) oled_data = 16'b0110101111000110;
    else if (pixel_index == 2173) oled_data = 16'b0101101101000010;
    else if (pixel_index == 2174) oled_data = 16'b0110110000000010;
    else if (pixel_index == 2175) oled_data = 16'b0101001111000001;
    else if (pixel_index == 2177 || pixel_index == 2278) oled_data = 16'b0100001100000010;
    else if (pixel_index == 2178) oled_data = 16'b0011001011000011;
    else if (pixel_index == 2180 || pixel_index == 3032) oled_data = 16'b0100001011000011;
    else if (pixel_index == 2181) oled_data = 16'b0011001010000000;
    else if (pixel_index == 2182) oled_data = 16'b0100101011000001;
    else if (pixel_index == 2185) oled_data = 16'b0110001111000011;
    else if (pixel_index == 2191) oled_data = 16'b0101001111000011;
    else if (pixel_index == 2192 || pixel_index == 2372) oled_data = 16'b0110010000000110;
    else if (pixel_index == 2196) oled_data = 16'b0011110010110110;
    else if (pixel_index == 2197 || ((pixel_index >= 2204) && (pixel_index <= 2207)) || pixel_index == 2228 || pixel_index == 2234 || pixel_index == 2316 || pixel_index == 2404 || pixel_index == 2594) oled_data = 16'b0011010010111011;
    else if (pixel_index == 2199 || ((pixel_index >= 2298) && (pixel_index <= 2299)) || pixel_index == 2302) oled_data = 16'b0011010011111100;
    else if (((pixel_index >= 2200) && (pixel_index <= 2201)) || pixel_index == 2505) oled_data = 16'b0010110011111100;
    else if (pixel_index == 2213) oled_data = 16'b0101110010110100;
    else if (pixel_index == 2214 || pixel_index == 2314) oled_data = 16'b0100110001010101;
    else if (pixel_index == 2215) oled_data = 16'b0100010001010101;
    else if (pixel_index == 2216 || pixel_index == 2604) oled_data = 16'b0101010001010100;
    else if (pixel_index == 2220) oled_data = 16'b0101110010110101;
    else if (pixel_index == 2224 || pixel_index == 2304 || pixel_index == 2313 || pixel_index == 3905) oled_data = 16'b0011110001011000;
    else if (pixel_index == 2226 || (pixel_index >= 2321) && (pixel_index <= 2322)) oled_data = 16'b0010010011111101;
    else if (pixel_index == 2227 || pixel_index == 2317) oled_data = 16'b0010010001011100;
    else if (pixel_index == 2230) oled_data = 16'b0001110010111110;
    else if (pixel_index == 2231) oled_data = 16'b0001110010111101;
    else if (pixel_index == 2233 || pixel_index == 2501) oled_data = 16'b0011010010111100;
    else if (pixel_index == 2236 || pixel_index == 2487) oled_data = 16'b0011110011111010;
    else if (pixel_index == 2237) oled_data = 16'b0100110011111010;
    else if (pixel_index == 2238) oled_data = 16'b0101110011110101;
    else if (pixel_index == 2242) oled_data = 16'b1000110100101110;
    else if (pixel_index == 2243) oled_data = 16'b1010010101101110;
    else if (pixel_index == 2246 || pixel_index == 2533 || pixel_index == 2815) oled_data = 16'b1000010100101110;
    else if (pixel_index == 2248 || pixel_index == 5329) oled_data = 16'b0111110000001111;
    else if (pixel_index == 2250 || pixel_index == 3461 || pixel_index == 4530) oled_data = 16'b0110101111010000;
    else if (pixel_index == 2251) oled_data = 16'b1000010000001101;
    else if (pixel_index == 2254) oled_data = 16'b0111101111001100;
    else if (pixel_index == 2256) oled_data = 16'b1001001111001011;
    else if (pixel_index == 2257 || pixel_index == 4750 || pixel_index == 5419) oled_data = 16'b1000001111001110;
    else if (pixel_index == 2258) oled_data = 16'b1001101111001101;
    else if (pixel_index == 2259) oled_data = 16'b0101001001000111;
    else if (pixel_index == 2260) oled_data = 16'b0110001010000110;
    else if (pixel_index == 2261) oled_data = 16'b0111101011001001;
    else if (pixel_index == 2262) oled_data = 16'b0110001101001100;
    else if (pixel_index == 2263 || pixel_index == 4176 || pixel_index == 4368) oled_data = 16'b0100001100001101;
    else if (pixel_index == 2266) oled_data = 16'b0111110001001100;
    else if (pixel_index == 2270) oled_data = 16'b0111110001000010;
    else if (pixel_index == 2271) oled_data = 16'b0110010001000011;
    else if (pixel_index == 2272) oled_data = 16'b0110010001000100;
    else if (pixel_index == 2273 || pixel_index == 2283) oled_data = 16'b0101101110000010;
    else if (pixel_index == 2274 || pixel_index == 2282) oled_data = 16'b0101001110000011;
    else if (pixel_index == 2275) oled_data = 16'b0101101111000110;
    else if (pixel_index == 2276 || pixel_index == 2676) oled_data = 16'b0101101101000100;
    else if (pixel_index == 2277) oled_data = 16'b0100001101000101;
    else if (pixel_index == 2280) oled_data = 16'b0101001110000100;
    else if (pixel_index == 2284 || pixel_index == 2381) oled_data = 16'b0101101111000100;
    else if (pixel_index == 2291) oled_data = 16'b0110110000001110;
    else if (pixel_index == 2292) oled_data = 16'b0110010001010011;
    else if (pixel_index == 2293 || pixel_index == 4003) oled_data = 16'b0100010001011000;
    else if (pixel_index == 2294 || pixel_index == 2323) oled_data = 16'b0011010010111010;
    else if (pixel_index == 2296 || pixel_index == 2410) oled_data = 16'b0010010100111011;
    else if (pixel_index == 2297) oled_data = 16'b0010110011111011;
    else if (((pixel_index >= 2300) && (pixel_index <= 2301)) || pixel_index == 2394 || ((pixel_index >= 2490) && (pixel_index <= 2491)) || pixel_index == 2493 || ((pixel_index >= 2587) && (pixel_index <= 2588)) || pixel_index == 2590 || pixel_index == 2687) oled_data = 16'b0011110100111100;
    else if (pixel_index == 2303 || pixel_index == 2393) oled_data = 16'b0011110011111100;
    else if (pixel_index == 2307) oled_data = 16'b0100110001010110;
    else if (pixel_index == 2308 || pixel_index == 3895) oled_data = 16'b0011110011111000;
    else if (pixel_index == 2309) oled_data = 16'b0100010100110111;
    else if (pixel_index == 2310) oled_data = 16'b0011010001011001;
    else if (pixel_index == 2311) oled_data = 16'b0011010000011010;
    else if (pixel_index == 2312) oled_data = 16'b0011010000011000;
    else if (pixel_index == 2319) oled_data = 16'b0001010010111011;
    else if (pixel_index == 2320) oled_data = 16'b0001010011111101;
    else if (pixel_index == 2324) oled_data = 16'b0010110010111001;
    else if (pixel_index == 2325 || pixel_index == 2593) oled_data = 16'b0011010010111001;
    else if (pixel_index == 2327) oled_data = 16'b0010110001010110;
    else if (pixel_index == 2328) oled_data = 16'b0010110010110101;
    else if (pixel_index == 2329 || pixel_index == 4320) oled_data = 16'b0100110011110101;
    else if (pixel_index == 2330) oled_data = 16'b0100110011110100;
    else if (pixel_index == 2331) oled_data = 16'b0100110011110010;
    else if (pixel_index == 2332) oled_data = 16'b0111010100101111;
    else if (pixel_index == 2333 || pixel_index == 2955) oled_data = 16'b1000010100101111;
    else if (pixel_index == 2334) oled_data = 16'b0110110011101000;
    else if (pixel_index == 2335 || pixel_index == 2426 || pixel_index == 2526 || pixel_index == 2991) oled_data = 16'b1000110011100111;
    else if (pixel_index == 2337) oled_data = 16'b1001010110100110;
    else if (pixel_index == 2338) oled_data = 16'b1010110110100111;
    else if (pixel_index == 2339 || pixel_index == 2529) oled_data = 16'b1010110110100110;
    else if (pixel_index == 2343) oled_data = 16'b0110010100110101;
    else if (pixel_index == 2344) oled_data = 16'b0101010001010101;
    else if (pixel_index == 2345 || pixel_index == 3817) oled_data = 16'b0101110011111000;
    else if (pixel_index == 2346) oled_data = 16'b0101110011110100;
    else if (pixel_index == 2347 || pixel_index == 2813 || pixel_index == 2969) oled_data = 16'b1000010100101101;
    else if (pixel_index == 2349) oled_data = 16'b1000110001000110;
    else if (pixel_index == 2350) oled_data = 16'b0111101101001001;
    else if (pixel_index == 2351) oled_data = 16'b0111101011001011;
    else if (pixel_index == 2352) oled_data = 16'b1000001011001010;
    else if (pixel_index == 2353) oled_data = 16'b0100100110000101;
    else if (pixel_index == 2354) oled_data = 16'b0110001000000110;
    else if (pixel_index == 2355 || pixel_index == 5326) oled_data = 16'b0110001001001001;
    else if (pixel_index == 2356) oled_data = 16'b0111001011001001;
    else if (pixel_index == 2357) oled_data = 16'b0110001011001001;
    else if (pixel_index == 2358) oled_data = 16'b0100101101001101;
    else if (pixel_index == 2360) oled_data = 16'b0011110001011010;
    else if (pixel_index == 2361 || pixel_index == 3835) oled_data = 16'b0101010100111010;
    else if (pixel_index == 2362 || pixel_index == 2855 || pixel_index == 2857 || pixel_index == 3221) oled_data = 16'b0111010110110111;
    else if (pixel_index == 2363) oled_data = 16'b0111110101110011;
    else if (pixel_index == 2368) oled_data = 16'b0111110011100111;
    else if (pixel_index == 2369 || pixel_index == 2616) oled_data = 16'b0111010000000011;
    else if (pixel_index == 2379) oled_data = 16'b0100001101000010;
    else if (pixel_index == 2380) oled_data = 16'b0101001110000101;
    else if (pixel_index == 2385) oled_data = 16'b0011001101001000;
    else if (pixel_index == 2387 || pixel_index == 2480) oled_data = 16'b0101110000001100;
    else if (pixel_index == 2390) oled_data = 16'b0100010010111011;
    else if (pixel_index == 2391) oled_data = 16'b0011110010111101;
    else if (pixel_index == 2392 || pixel_index == 2506) oled_data = 16'b0011010011111101;
    else if (((pixel_index >= 2395) && (pixel_index <= 2396)) || ((pixel_index >= 2398) && (pixel_index <= 2399)) || pixel_index == 2411 || pixel_index == 2492 || pixel_index == 2502) oled_data = 16'b0011010100111100;
    else if (pixel_index == 2397 || pixel_index == 2507) oled_data = 16'b0011110100111101;
    else if (pixel_index == 2401) oled_data = 16'b0010001111010100;
    else if (pixel_index == 2402) oled_data = 16'b0010110001011000;
    else if (pixel_index == 2403) oled_data = 16'b0011110010111010;
    else if (pixel_index == 2405) oled_data = 16'b0011010011111010;
    else if (pixel_index == 2409) oled_data = 16'b0010110010111101;
    else if (pixel_index == 2412) oled_data = 16'b0010110100111100;
    else if (pixel_index == 2413 || pixel_index == 3891 || pixel_index == 3957) oled_data = 16'b0010110100111010;
    else if ((pixel_index >= 2414) && (pixel_index <= 2415)) oled_data = 16'b0010110011111010;
    else if (pixel_index == 2417 || pixel_index == 2757) oled_data = 16'b0110110100110101;
    else if (pixel_index == 2419 || pixel_index == 2776) oled_data = 16'b0110110001001101;
    else if (pixel_index == 2429 || pixel_index == 2805) oled_data = 16'b0111110011100101;
    else if (pixel_index == 2430) oled_data = 16'b0111110011100011;
    else if (pixel_index == 2431) oled_data = 16'b1000110011100011;
    else if (pixel_index == 2434 || pixel_index == 3086) oled_data = 16'b1010010110101011;
    else if (pixel_index == 2435 || pixel_index == 3090) oled_data = 16'b1001010111101001;
    else if (pixel_index == 2438 || pixel_index == 2460) oled_data = 16'b0110110100110001;
    else if (pixel_index == 2440 || pixel_index == 2826 || pixel_index == 2829) oled_data = 16'b0101010001010000;
    else if (pixel_index == 2441 || pixel_index == 3059) oled_data = 16'b0110110011110000;
    else if (pixel_index == 2443) oled_data = 16'b1010010100101010;
    else if (pixel_index == 2444) oled_data = 16'b1001110010101000;
    else if (pixel_index == 2445) oled_data = 16'b0111001110000100;
    else if (pixel_index == 2446) oled_data = 16'b0110001011000110;
    else if (pixel_index == 2447) oled_data = 16'b0101100111000101;
    else if (pixel_index == 2448 || pixel_index == 2646) oled_data = 16'b0101000110000100;
    else if (pixel_index == 2449) oled_data = 16'b0100100101000011;
    else if (pixel_index == 2450) oled_data = 16'b0100100101000100;
    else if (pixel_index == 2451) oled_data = 16'b0100000100000011;
    else if (pixel_index == 2452) oled_data = 16'b0100000110000100;
    else if (pixel_index == 2453 || pixel_index == 2542 || pixel_index == 2746) oled_data = 16'b0100101000000101;
    else if (pixel_index == 2454) oled_data = 16'b0101101011001001;
    else if (pixel_index == 2455) oled_data = 16'b0101001111010100;
    else if (pixel_index == 2456 || pixel_index == 3906) oled_data = 16'b0011110001011001;
    else if (pixel_index == 2457 || pixel_index == 2586 || (pixel_index >= 2684) && (pixel_index <= 2685)) oled_data = 16'b0100010101111101;
    else if (pixel_index == 2458) oled_data = 16'b0101010101111110;
    else if (pixel_index == 2459) oled_data = 16'b0111010101110110;
    else if (pixel_index == 2461 || pixel_index == 2628) oled_data = 16'b0111110011101100;
    else if (pixel_index == 2462) oled_data = 16'b0111110010101100;
    else if (pixel_index == 2468 || pixel_index == 2471) oled_data = 16'b0110010000001000;
    else if (pixel_index == 2469 || pixel_index == 2472) oled_data = 16'b0101010000001010;
    else if (pixel_index == 2479) oled_data = 16'b0101001110001000;
    else if (pixel_index == 2482) oled_data = 16'b0011101110000111;
    else if (pixel_index == 2485) oled_data = 16'b0011110001010010;
    else if (pixel_index == 2486) oled_data = 16'b0011110011110101;
    else if (pixel_index == 2488 || pixel_index == 2690) oled_data = 16'b0011110100111011;
    else if (pixel_index == 2489 || pixel_index == 2686) oled_data = 16'b0011110101111100;
    else if (pixel_index == 2494 || pixel_index == 2683 || pixel_index == 2696) oled_data = 16'b0100010100111101;
    else if (pixel_index == 2495 || pixel_index == 2589) oled_data = 16'b0100010100111100;
    else if (pixel_index == 2499) oled_data = 16'b0011110001010011;
    else if (pixel_index == 2500) oled_data = 16'b0100010001011001;
    else if ((pixel_index >= 2503) && (pixel_index <= 2504)) oled_data = 16'b0010110101111100;
    else if (pixel_index == 2508 || pixel_index == 2681) oled_data = 16'b0100110100111001;
    else if (pixel_index == 2509 || pixel_index == 4092) oled_data = 16'b0101010100110100;
    else if (pixel_index == 2511) oled_data = 16'b0111010001001101;
    else if (pixel_index == 2513 || pixel_index == 3082) oled_data = 16'b1010010011101010;
    else if (pixel_index == 2514) oled_data = 16'b1001110011101001;
    else if (pixel_index == 2520) oled_data = 16'b1001110100100100;
    else if (pixel_index == 2523) oled_data = 16'b1001010011100100;
    else if (pixel_index == 2527) oled_data = 16'b1000110011100100;
    else if (pixel_index == 2530) oled_data = 16'b1001010101100100;
    else if (pixel_index == 2531) oled_data = 16'b0111110101101001;
    else if (pixel_index == 2532) oled_data = 16'b0111010100101100;
    else if (pixel_index == 2534 || pixel_index == 2796) oled_data = 16'b0111110011101110;
    else if (pixel_index == 2536 || pixel_index == 2540) oled_data = 16'b0101101100000111;
    else if (pixel_index == 2537) oled_data = 16'b0110001101000101;
    else if (pixel_index == 2538) oled_data = 16'b0110001011000011;
    else if (pixel_index == 2539 || pixel_index == 3230) oled_data = 16'b0110001100000111;
    else if (pixel_index == 2541 || pixel_index == 2642) oled_data = 16'b0100000111000100;
    else if (pixel_index == 2543) oled_data = 16'b0100100110000100;
    else if (pixel_index == 2544 || pixel_index == 3172 || pixel_index == 3696 || pixel_index == 3983) oled_data = 16'b0011000110000101;
    else if (pixel_index == 2545) oled_data = 16'b0100000110000101;
    else if (pixel_index == 2546 || pixel_index == 3600 || pixel_index == 3887) oled_data = 16'b0010100100000011;
    else if (pixel_index == 2547) oled_data = 16'b0011000011000001;
    else if (pixel_index == 2548) oled_data = 16'b0011000011000011;
    else if (pixel_index == 2549) oled_data = 16'b0100100111000011;
    else if (pixel_index == 2550) oled_data = 16'b0111101010000101;
    else if (pixel_index == 2551) oled_data = 16'b1010101110001000;
    else if (pixel_index == 2552) oled_data = 16'b1000101110001011;
    else if (pixel_index == 2554 || pixel_index == 2694) oled_data = 16'b0100110100111010;
    else if (pixel_index == 2555) oled_data = 16'b0101110101111100;
    else if (pixel_index == 2556) oled_data = 16'b0110010100110111;
    else if (pixel_index == 2557) oled_data = 16'b0111010100110001;
    else if (pixel_index == 2558) oled_data = 16'b0111110100110100;
    else if (pixel_index == 2560 || pixel_index == 3096) oled_data = 16'b1000010011101110;
    else if (pixel_index == 2562) oled_data = 16'b0110010001001110;
    else if (pixel_index == 2565 || pixel_index == 2664) oled_data = 16'b0100110000010000;
    else if (pixel_index == 2568) oled_data = 16'b0100110000001101;
    else if (pixel_index == 2571) oled_data = 16'b0101101101000011;
    else if (pixel_index == 2575) oled_data = 16'b0100101111000110;
    else if (pixel_index == 2577 || pixel_index == 3420) oled_data = 16'b0110110010101101;
    else if (pixel_index == 2578) oled_data = 16'b0101101111001001;
    else if (pixel_index == 2582) oled_data = 16'b0100110001001101;
    else if (pixel_index == 2583) oled_data = 16'b0101010011110011;
    else if (pixel_index == 2584) oled_data = 16'b0100110101111010;
    else if (pixel_index == 2585) oled_data = 16'b0100110100111101;
    else if (pixel_index == 2591) oled_data = 16'b0100010011111100;
    else if (pixel_index == 2595) oled_data = 16'b0010110100111011;
    else if (pixel_index == 2596) oled_data = 16'b0011010101111101;
    else if ((pixel_index >= 2597) && (pixel_index <= 2598)) oled_data = 16'b0011010100111101;
    else if ((pixel_index >= 2599) && (pixel_index <= 2600)) oled_data = 16'b0010110110111101;
    else if (pixel_index == 2601 || pixel_index == 2692) oled_data = 16'b0011010101111100;
    else if (pixel_index == 2602) oled_data = 16'b0100010100111011;
    else if (pixel_index == 2603 || pixel_index == 3999) oled_data = 16'b0100110011111000;
    else if (pixel_index == 2606) oled_data = 16'b0101101101001011;
    else if (pixel_index == 2607) oled_data = 16'b0110101110001001;
    else if (pixel_index == 2608) oled_data = 16'b1000110000000111;
    else if (pixel_index == 2609) oled_data = 16'b1000001111000101;
    else if (pixel_index == 2614 || pixel_index == 2623) oled_data = 16'b1001110101100110;
    else if (pixel_index == 2621) oled_data = 16'b1001010101101001;
    else if (pixel_index == 2622 || pixel_index == 3055) oled_data = 16'b1000110011101010;
    else if (pixel_index == 2624) oled_data = 16'b1001110110101000;
    else if (pixel_index == 2627) oled_data = 16'b0110110101101101;
    else if (pixel_index == 2631 || pixel_index == 2726) oled_data = 16'b0110101101000111;
    else if (pixel_index == 2632 || pixel_index == 2728 || pixel_index == 2745) oled_data = 16'b0100001001000010;
    else if (pixel_index == 2633) oled_data = 16'b0100001001000000;
    else if (pixel_index == 2634) oled_data = 16'b0011101000000001;
    else if (pixel_index == 2635) oled_data = 16'b0010100111000100;
    else if (pixel_index == 2636) oled_data = 16'b0010100110000100;
    else if (pixel_index == 2637) oled_data = 16'b0011100101000011;
    else if (pixel_index == 2638) oled_data = 16'b0101101010000111;
    else if (pixel_index == 2640) oled_data = 16'b0101101010001000;
    else if (pixel_index == 2641) oled_data = 16'b0100100111000101;
    else if (pixel_index == 2643) oled_data = 16'b0101001000000101;
    else if (pixel_index == 2644) oled_data = 16'b0110001001000110;
    else if (pixel_index == 2645 || pixel_index == 2833) oled_data = 16'b0101000111000111;
    else if (pixel_index == 2647) oled_data = 16'b0111101010000011;
    else if (pixel_index == 2648) oled_data = 16'b1000001101000100;
    else if (pixel_index == 2649 || pixel_index == 2736) oled_data = 16'b0110001010001000;
    else if (pixel_index == 2650) oled_data = 16'b0100001111010010;
    else if (pixel_index == 2651 || pixel_index == 3825 || pixel_index == 3831) oled_data = 16'b0101010100111011;
    else if (pixel_index == 2652 || pixel_index == 3753) oled_data = 16'b0101110101111011;
    else if (pixel_index == 2653 || pixel_index == 3007 || pixel_index == 3220) oled_data = 16'b0111110111111011;
    else if (pixel_index == 2654 || pixel_index == 2920 || pixel_index == 3771 || pixel_index == 3799) oled_data = 16'b0110010110111011;
    else if (pixel_index == 2655) oled_data = 16'b0111010100110111;
    else if (pixel_index == 2656) oled_data = 16'b1001010100110010;
    else if (pixel_index == 2657) oled_data = 16'b1000110100101111;
    else if (pixel_index == 2659) oled_data = 16'b0110010110111000;
    else if (pixel_index == 2660) oled_data = 16'b0110010010110001;
    else if (pixel_index == 2662) oled_data = 16'b0101001111001110;
    else if (pixel_index == 2666) oled_data = 16'b0101001110001010;
    else if (pixel_index == 2667) oled_data = 16'b0101101011000011;
    else if (pixel_index == 2673) oled_data = 16'b0110010010101101;
    else if (pixel_index == 2678) oled_data = 16'b0101101110000110;
    else if (pixel_index == 2680 || pixel_index == 2777) oled_data = 16'b0110010011110011;
    else if (pixel_index == 2682) oled_data = 16'b0100010101111100;
    else if (pixel_index == 2689) oled_data = 16'b0011010101111011;
    else if (pixel_index == 2691) oled_data = 16'b0100010101111110;
    else if (pixel_index == 2693) oled_data = 16'b0100110101111011;
    else if (pixel_index == 2695) oled_data = 16'b0100110101111101;
    else if (pixel_index == 2697) oled_data = 16'b0100010011111010;
    else if (pixel_index == 2698) oled_data = 16'b0101110100111000;
    else if (pixel_index == 2700) oled_data = 16'b0110001111001110;
    else if (pixel_index == 2701) oled_data = 16'b0111001111001011;
    else if (pixel_index == 2703) oled_data = 16'b1000010000001011;
    else if (pixel_index == 2704) oled_data = 16'b1000010001001010;
    else if (pixel_index == 2712) oled_data = 16'b0111010001000011;
    else if (pixel_index == 2714) oled_data = 16'b1000010011100100;
    else if (pixel_index == 2715 || pixel_index == 2807) oled_data = 16'b0111010010100011;
    else if (pixel_index == 2719) oled_data = 16'b1000110101101011;
    else if (pixel_index == 2720) oled_data = 16'b1000110100101100;
    else if (pixel_index == 2727) oled_data = 16'b0101101010000011;
    else if (pixel_index == 2729) oled_data = 16'b0011101000000010;
    else if (pixel_index == 2732) oled_data = 16'b0010000101000100;
    else if (pixel_index == 2733) oled_data = 16'b0100001001000011;
    else if (pixel_index == 2735) oled_data = 16'b0110101110001101;
    else if (pixel_index == 2737 || pixel_index == 3268) oled_data = 16'b0011000111000111;
    else if (pixel_index == 2738) oled_data = 16'b0101000110001000;
    else if (pixel_index == 2739 || pixel_index == 2840) oled_data = 16'b1001001110001100;
    else if (pixel_index == 2740) oled_data = 16'b1001101110001011;
    else if (pixel_index == 2741) oled_data = 16'b1000001101001010;
    else if (pixel_index == 2742) oled_data = 16'b0101000111000101;
    else if (pixel_index == 2743) oled_data = 16'b0100100110000011;
    else if (pixel_index == 2744) oled_data = 16'b0101001010000101;
    else if (pixel_index == 2747 || pixel_index == 2825) oled_data = 16'b0101001111001111;
    else if (pixel_index == 2748 || pixel_index == 3987) oled_data = 16'b0110010101111010;
    else if (pixel_index == 2749) oled_data = 16'b0110010110111110;
    else if (pixel_index == 2750 || pixel_index == 2779) oled_data = 16'b0101010101111101;
    else if (pixel_index == 2751 || pixel_index == 3788) oled_data = 16'b0101110111111011;
    else if (pixel_index == 2752) oled_data = 16'b1000010110111001;
    else if (pixel_index == 2753) oled_data = 16'b0111110101111010;
    else if (pixel_index == 2754 || pixel_index == 2793 || pixel_index == 3757 || pixel_index == 3779 || pixel_index == 3784 || pixel_index == 3797) oled_data = 16'b0110010110111010;
    else if (pixel_index == 2755 || pixel_index == 3782) oled_data = 16'b0110110111111011;
    else if (pixel_index == 2756) oled_data = 16'b0111110100110110;
    else if (pixel_index == 2758) oled_data = 16'b0110110010110011;
    else if (pixel_index == 2759 || pixel_index == 2761 || pixel_index == 4089) oled_data = 16'b0110110100110011;
    else if (pixel_index == 2760 || pixel_index == 2917) oled_data = 16'b0110010100110011;
    else if (pixel_index == 2762 || pixel_index == 3058) oled_data = 16'b0110010001001101;
    else if (pixel_index == 2763) oled_data = 16'b0101101100000100;
    else if (pixel_index == 2765) oled_data = 16'b0101110010101101;
    else if (pixel_index == 2774 || pixel_index == 3093) oled_data = 16'b0110101110000011;
    else if (pixel_index == 2778 || pixel_index == 2792 || pixel_index == 3823 || pixel_index == 3978) oled_data = 16'b0101010101111011;
    else if (pixel_index == 2780) oled_data = 16'b0101010110111100;
    else if (pixel_index == 2781 || pixel_index == 3795) oled_data = 16'b0101010101111100;
    else if (pixel_index == 2782) oled_data = 16'b0101010110111101;
    else if (pixel_index == 2783) oled_data = 16'b0100110101111100;
    else if (pixel_index == 2784) oled_data = 16'b0010001111010101;
    else if (pixel_index == 2785 || pixel_index == 3879 || pixel_index == 3893) oled_data = 16'b0010110011111001;
    else if (pixel_index == 2789) oled_data = 16'b0101010011110110;
    else if (pixel_index == 2790 || pixel_index == 3812 || pixel_index == 3814 || pixel_index == 3816) oled_data = 16'b0101010011111000;
    else if (pixel_index == 2791 || pixel_index == 2845) oled_data = 16'b0101010101111010;
    else if (pixel_index == 2794) oled_data = 16'b0111110110110110;
    else if (pixel_index == 2795) oled_data = 16'b1001010110110010;
    else if (pixel_index == 2798) oled_data = 16'b0110110001001011;
    else if (pixel_index == 2802) oled_data = 16'b1001010011101011;
    else if (pixel_index == 2804) oled_data = 16'b0111010010100101;
    else if (pixel_index == 2806) oled_data = 16'b0111110100100101;
    else if (pixel_index == 2814) oled_data = 16'b0111110100101110;
    else if (pixel_index == 2816) oled_data = 16'b1000010101101111;
    else if (pixel_index == 2818 || pixel_index == 3154) oled_data = 16'b1000010001001101;
    else if (pixel_index == 2827) oled_data = 16'b0101110000010000;
    else if (pixel_index == 2828) oled_data = 16'b0101001110001110;
    else if (pixel_index == 2830) oled_data = 16'b0101110100110110;
    else if (pixel_index == 2831) oled_data = 16'b0110110010110101;
    else if (pixel_index == 2832) oled_data = 16'b0101001001001011;
    else if (pixel_index == 2834) oled_data = 16'b0101100111000110;
    else if (pixel_index == 2835) oled_data = 16'b1000101100001000;
    else if (pixel_index == 2836) oled_data = 16'b0111101100000111;
    else if (pixel_index == 2837) oled_data = 16'b0111001011000110;
    else if (pixel_index == 2838) oled_data = 16'b1000001000000100;
    else if (pixel_index == 2839) oled_data = 16'b1001001100001001;
    else if (pixel_index == 2841) oled_data = 16'b0101001001000100;
    else if (pixel_index == 2842) oled_data = 16'b0011100110000001;
    else if (pixel_index == 2846 || pixel_index == 3019) oled_data = 16'b0110010111111101;
    else if (pixel_index == 2847 || pixel_index == 3018) oled_data = 16'b0101111000111110;
    else if (pixel_index == 2848 || pixel_index == 3014) oled_data = 16'b0110110110111101;
    else if (pixel_index == 2849) oled_data = 16'b0111010111111111;
    else if (pixel_index == 2850) oled_data = 16'b0110010111111111;
    else if (pixel_index == 2851 || pixel_index == 3115) oled_data = 16'b0110110111111101;
    else if (pixel_index == 2852 || pixel_index == 2952 || pixel_index == 3100) oled_data = 16'b0111110110111010;
    else if (pixel_index == 2853) oled_data = 16'b0111010110111001;
    else if (pixel_index == 2854) oled_data = 16'b0111010101111000;
    else if (pixel_index == 2856 || pixel_index == 3005) oled_data = 16'b0111110101110101;
    else if (pixel_index == 2859) oled_data = 16'b0111001111000111;
    else if (pixel_index == 2873 || pixel_index == 3105) oled_data = 16'b0111110100110000;
    else if (pixel_index == 2874 || pixel_index == 3038) oled_data = 16'b0110110101111000;
    else if (pixel_index == 2875 || ((pixel_index >= 2877) && (pixel_index <= 2878)) || pixel_index == 3763) oled_data = 16'b0101110110111100;
    else if (pixel_index == 2876) oled_data = 16'b0101110110111101;
    else if (pixel_index == 2879) oled_data = 16'b0101110111111101;
    else if (pixel_index == 2880 || pixel_index == 5988) oled_data = 16'b0011001001001011;
    else if (pixel_index == 2884) oled_data = 16'b0100110000010011;
    else if (pixel_index == 2885) oled_data = 16'b0100010011110110;
    else if (pixel_index == 2886) oled_data = 16'b0101010100110111;
    else if (pixel_index == 2887) oled_data = 16'b0100110100110101;
    else if (pixel_index == 2889 || pixel_index == 3750) oled_data = 16'b0101110100110111;
    else if (pixel_index == 2891) oled_data = 16'b1000010100110011;
    else if (pixel_index == 2892) oled_data = 16'b1000010010110001;
    else if (pixel_index == 2893) oled_data = 16'b0110110001001111;
    else if (pixel_index == 2898) oled_data = 16'b1001110110101001;
    else if (pixel_index == 2900) oled_data = 16'b0111010000000001;
    else if (pixel_index == 2902) oled_data = 16'b0110110011100011;
    else if (pixel_index == 2903) oled_data = 16'b0110110010100110;
    else if (pixel_index == 2909 || pixel_index == 3708) oled_data = 16'b1000110101110010;
    else if (pixel_index == 2910) oled_data = 16'b1000010101110011;
    else if (pixel_index == 2911) oled_data = 16'b1000010101110010;
    else if (pixel_index == 2912 || pixel_index == 5364) oled_data = 16'b1001010110110101;
    else if (pixel_index == 2913) oled_data = 16'b1001010110110000;
    else if (pixel_index == 2914) oled_data = 16'b1001010000001001;
    else if (pixel_index == 2915) oled_data = 16'b0110101110000111;
    else if (pixel_index == 2921) oled_data = 16'b0101010111111101;
    else if (pixel_index == 2922 || pixel_index == 2926) oled_data = 16'b0110111000111111;
    else if (pixel_index == 2923 || pixel_index == 3020 || (pixel_index >= 3109) && (pixel_index <= 3110)) oled_data = 16'b0110111000111110;
    else if (pixel_index == 2924 || pixel_index == 2945 || pixel_index == 3040 || pixel_index == 3103) oled_data = 16'b0111011000111100;
    else if (pixel_index == 2925) oled_data = 16'b0101110111111111;
    else if (pixel_index == 2927) oled_data = 16'b0110110101110110;
    else if (pixel_index == 2928 || pixel_index == 4079) oled_data = 16'b0100000111000111;
    else if (pixel_index == 2929) oled_data = 16'b0100100100000101;
    else if (pixel_index == 2931) oled_data = 16'b1001001111001010;
    else if (pixel_index == 2932) oled_data = 16'b0110100111000100;
    else if (pixel_index == 2933) oled_data = 16'b0101100110000100;
    else if (pixel_index == 2934 || pixel_index == 3029) oled_data = 16'b1001101101001000;
    else if (pixel_index == 2935) oled_data = 16'b1010110000001010;
    else if (pixel_index == 2936 || pixel_index == 3273) oled_data = 16'b1000001110001001;
    else if (pixel_index == 2937) oled_data = 16'b0011000111000010;
    else if (pixel_index == 2938) oled_data = 16'b0001000111000001;
    else if (pixel_index == 2939) oled_data = 16'b0011001000000011;
    else if (pixel_index == 2941) oled_data = 16'b0100101111010011;
    else if (pixel_index == 2942) oled_data = 16'b0110111000111101;
    else if (pixel_index == 2943 || pixel_index == 3016 || pixel_index == 3022) oled_data = 16'b0111011000111110;
    else if (pixel_index == 2944 || pixel_index == 3071) oled_data = 16'b0111010111111100;
    else if (pixel_index == 2946) oled_data = 16'b0110011000111101;
    else if (pixel_index == 2947) oled_data = 16'b0110110111111110;
    else if (pixel_index == 2948 || pixel_index == 3015 || pixel_index == 3017 || pixel_index == 3111) oled_data = 16'b0110010111111110;
    else if (pixel_index == 2949 || pixel_index == 3102) oled_data = 16'b0111010111111110;
    else if (pixel_index == 2950 || pixel_index == 3069) oled_data = 16'b0111010111111101;
    else if (pixel_index == 2951 || pixel_index == 3070) oled_data = 16'b0111110111111100;
    else if (pixel_index == 2953) oled_data = 16'b1000010110111100;
    else if (pixel_index == 2954) oled_data = 16'b0111010100110101;
    else if (pixel_index == 2956) oled_data = 16'b1000110101110001;
    else if (pixel_index == 2957 || pixel_index == 3155 || pixel_index == 3462) oled_data = 16'b0111110011110001;
    else if (pixel_index == 2970) oled_data = 16'b0111010100110100;
    else if (pixel_index == 2971 || pixel_index == 3770) oled_data = 16'b0110110110111010;
    else if (pixel_index == 2972 || pixel_index == 2974 || pixel_index == 3101 || pixel_index == 3986) oled_data = 16'b0110110110111011;
    else if (pixel_index == 2973 || pixel_index == 3042 || ((pixel_index >= 3767) && (pixel_index <= 3768)) || pixel_index == 3781 || pixel_index == 4471) oled_data = 16'b0110110111111100;
    else if (pixel_index == 2975 || pixel_index == 3107) oled_data = 16'b0111010110111011;
    else if (pixel_index == 2976) oled_data = 16'b0011001010001011;
    else if (pixel_index == 2978) oled_data = 16'b0100101101001111;
    else if (pixel_index == 2981 || pixel_index == 3778) oled_data = 16'b0110110110111000;
    else if (pixel_index == 2982 || pixel_index == 4184 || pixel_index == 4460) oled_data = 16'b0111010111111001;
    else if (pixel_index == 2983 || pixel_index == 3657) oled_data = 16'b1000010100110100;
    else if (pixel_index == 2985) oled_data = 16'b0111010000001110;
    else if (pixel_index == 2986) oled_data = 16'b1000110001001010;
    else if (pixel_index == 2987) oled_data = 16'b1001010001001001;
    else if (pixel_index == 2988) oled_data = 16'b1000010000001010;
    else if (pixel_index == 2990) oled_data = 16'b1000010010101011;
    else if (pixel_index == 2992) oled_data = 16'b1000010101101010;
    else if (pixel_index == 2993) oled_data = 16'b1000010110101011;
    else if (pixel_index == 2994) oled_data = 16'b1000110110100110;
    else if (pixel_index == 2997) oled_data = 16'b0110001110000000;
    else if (pixel_index == 2998) oled_data = 16'b0110110001000110;
    else if (pixel_index == 3004) oled_data = 16'b0111110110110011;
    else if (pixel_index == 3006) oled_data = 16'b0111010111111010;
    else if (pixel_index == 3008 || pixel_index == 4447) oled_data = 16'b1000010111111011;
    else if (pixel_index == 3009) oled_data = 16'b1000010101110000;
    else if (pixel_index == 3010) oled_data = 16'b0111110000001001;
    else if (pixel_index == 3011) oled_data = 16'b0111010011110101;
    else if (pixel_index == 3012) oled_data = 16'b0110110101111011;
    else if (pixel_index == 3013) oled_data = 16'b0110110110111111;
    else if (pixel_index == 3021 || pixel_index == 3116 || pixel_index == 3776) oled_data = 16'b0111011001111110;
    else if (pixel_index == 3023) oled_data = 16'b0110110001010110;
    else if (pixel_index == 3027) oled_data = 16'b1001010110111010;
    else if (pixel_index == 3028) oled_data = 16'b1000101110001101;
    else if (pixel_index == 3030) oled_data = 16'b1001110000001101;
    else if (pixel_index == 3031) oled_data = 16'b0110101100001001;
    else if (pixel_index == 3033) oled_data = 16'b0010100111000000;
    else if (pixel_index == 3034) oled_data = 16'b0010000110000000;
    else if (pixel_index == 3035) oled_data = 16'b0011100111000110;
    else if (pixel_index == 3039) oled_data = 16'b0111111001111110;
    else if (pixel_index == 3041 || pixel_index == 4472 || pixel_index == 4477 || pixel_index == 4488) oled_data = 16'b0110111000111100;
    else if (pixel_index == 3043 || pixel_index == 3775) oled_data = 16'b0111011000111011;
    else if (pixel_index == 3044 || pixel_index == 3139 || pixel_index == 4582) oled_data = 16'b1001011000111100;
    else if (pixel_index == 3045 || pixel_index == 3509 || pixel_index == 3578 || pixel_index == 3596 || pixel_index == 3688 || pixel_index == 3702) oled_data = 16'b1010011010111110;
    else if (pixel_index == 3046 || pixel_index == 3234 || pixel_index == 3497 || pixel_index == 3507 || pixel_index == 3534 || pixel_index == 3603 || pixel_index == 3620 || pixel_index == 3674 || pixel_index == 3678 || pixel_index == 3691) oled_data = 16'b1010111001111101;
    else if (pixel_index == 3047 || pixel_index == 3147 || pixel_index == 3243 || pixel_index == 3262 || pixel_index == 3359 || pixel_index == 3402 || (pixel_index >= 3435) && (pixel_index <= 3437)) oled_data = 16'b1011111010111101;
    else if (pixel_index == 3048 || pixel_index == 3244 || pixel_index == 3335 || pixel_index == 3338 || pixel_index == 3355 || pixel_index == 3357 || pixel_index == 3393 || pixel_index == 3431 || pixel_index == 4696) oled_data = 16'b1100011011111101;
    else if (pixel_index == 3049 || pixel_index == 3439 || pixel_index == 4566) oled_data = 16'b1010111010111011;
    else if (pixel_index == 3050) oled_data = 16'b1010011000111011;
    else if (pixel_index == 3051) oled_data = 16'b1001110111111001;
    else if (pixel_index == 3052) oled_data = 16'b1001111000111001;
    else if (pixel_index == 3053) oled_data = 16'b1000110100110101;
    else if (pixel_index == 3060) oled_data = 16'b0110010000001011;
    else if (pixel_index == 3066 || pixel_index == 3561 || pixel_index == 3711) oled_data = 16'b1000010101110101;
    else if (pixel_index == 3067) oled_data = 16'b0111110110111011;
    else if (pixel_index == 3068) oled_data = 16'b0111110111111101;
    else if (pixel_index == 3074) oled_data = 16'b0100010011110111;
    else if (pixel_index == 3075) oled_data = 16'b0100010101110111;
    else if (pixel_index == 3076) oled_data = 16'b0100110011110111;
    else if (pixel_index == 3077) oled_data = 16'b0111111000111010;
    else if (pixel_index == 3078 || pixel_index == 3164 || pixel_index == 3545 || pixel_index == 3549 || ((pixel_index >= 3569) && (pixel_index <= 3570)) || pixel_index == 3572 || pixel_index == 3633 || pixel_index == 3667 || ((pixel_index >= 3737) && (pixel_index <= 3738)) || pixel_index == 4602) oled_data = 16'b1001111010111101;
    else if (pixel_index == 3079) oled_data = 16'b1010011000111001;
    else if (pixel_index == 3081) oled_data = 16'b1000110001001100;
    else if (pixel_index == 3083) oled_data = 16'b1010010011101001;
    else if (pixel_index == 3084) oled_data = 16'b1010010010101011;
    else if (pixel_index == 3085) oled_data = 16'b1010010101101100;
    else if (pixel_index == 3087) oled_data = 16'b1010010111101010;
    else if (pixel_index == 3088) oled_data = 16'b1010010111101101;
    else if (pixel_index == 3089) oled_data = 16'b1001010111101101;
    else if (pixel_index == 3094) oled_data = 16'b1000001111000111;
    else if (pixel_index == 3097 || pixel_index == 3517) oled_data = 16'b0111110001001111;
    else if (pixel_index == 3099) oled_data = 16'b1000110100110100;
    else if (pixel_index == 3104) oled_data = 16'b0111010111111000;
    else if (pixel_index == 3108 || pixel_index == 3112 || pixel_index == 4476) oled_data = 16'b0111011000111101;
    else if (pixel_index == 3113) oled_data = 16'b1000010111111101;
    else if (pixel_index == 3114 || pixel_index == 4450) oled_data = 16'b0111111000111100;
    else if (pixel_index == 3117) oled_data = 16'b0111111000111110;
    else if (pixel_index == 3118 || pixel_index == 3138 || pixel_index == 3495 || pixel_index == 3548 || pixel_index == 3551 || pixel_index == 3568 || pixel_index == 3584 || pixel_index == 3619 || pixel_index == 3714) oled_data = 16'b1010011001111100;
    else if (pixel_index == 3120) oled_data = 16'b0100100110000110;
    else if (pixel_index == 3121 || pixel_index == 3792) oled_data = 16'b0010100101000100;
    else if (pixel_index == 3122) oled_data = 16'b0110110010110110;
    else if (pixel_index == 3123) oled_data = 16'b0111011001111111;
    else if (pixel_index == 3124) oled_data = 16'b0111010001010011;
    else if (pixel_index == 3125) oled_data = 16'b1000110010110001;
    else if (pixel_index == 3127 || pixel_index == 3557) oled_data = 16'b0101101100001011;
    else if (pixel_index == 3128) oled_data = 16'b0011001001000100;
    else if (pixel_index == 3130) oled_data = 16'b0010000110000010;
    else if (pixel_index == 3131) oled_data = 16'b0011100111000001;
    else if (pixel_index == 3132) oled_data = 16'b0101001001000011;
    else if (pixel_index == 3133) oled_data = 16'b0101001011000111;
    else if (pixel_index == 3135 || pixel_index == 3426 || pixel_index == 3449 || pixel_index == 3455 || pixel_index == 3523 || pixel_index == 3533 || pixel_index == 3565 || pixel_index == 3594 || pixel_index == 3685 || pixel_index == 3692 || pixel_index == 3715 || pixel_index == 4569) oled_data = 16'b1010111010111100;
    else if (pixel_index == 3136 || pixel_index == 3219 || pixel_index == 3477 || pixel_index == 3573 || pixel_index == 3662 || ((pixel_index >= 3668) && (pixel_index <= 3669)) || pixel_index == 3722 || pixel_index == 3735) oled_data = 16'b1001111010111110;
    else if (pixel_index == 3137 || pixel_index == 3739) oled_data = 16'b1001011001111110;
    else if (pixel_index == 3140 || pixel_index == 3680 || pixel_index == 4568) oled_data = 16'b1011011011111100;
    else if (pixel_index == 3141 || pixel_index == 3308 || pixel_index == 4548 || pixel_index == 4673 || ((pixel_index >= 4687) && (pixel_index <= 4689)) || pixel_index == 5188 || pixel_index == 5478) oled_data = 16'b1101011100111100;
    else if (pixel_index == 3142 || pixel_index == 4664 || pixel_index == 4679 || pixel_index == 4681 || pixel_index == 4807 || pixel_index == 4894 || pixel_index == 4957 || pixel_index == 4963 || pixel_index == 5009 || pixel_index == 5123 || pixel_index == 5380 || pixel_index == 5614 || pixel_index == 6121) oled_data = 16'b1101111100111101;
    else if (pixel_index == 3143 || pixel_index == 4662 || pixel_index == 5187 || pixel_index == 5197 || pixel_index == 5288 || pixel_index == 5394 || ((pixel_index >= 5523) && (pixel_index <= 5524)) || pixel_index == 5581 || pixel_index == 5597 || pixel_index == 5700 || (pixel_index >= 5773) && (pixel_index <= 5774)) oled_data = 16'b1110011101111100;
    else if (pixel_index == 3144 || pixel_index == 4745 || pixel_index == 4782 || pixel_index == 4843 || pixel_index == 5097 || pixel_index == 5294 || pixel_index == 5302 || pixel_index == 5308 || pixel_index == 5389 || pixel_index == 5400 || pixel_index == 5491 || pixel_index == 5549 || pixel_index == 5593 || pixel_index == 5725 || pixel_index == 5820 || pixel_index == 6020) oled_data = 16'b1110111110111101;
    else if (pixel_index == 3145) oled_data = 16'b1100111101111101;
    else if (pixel_index == 3146 || pixel_index == 3290 || pixel_index == 3332 || pixel_index == 3412) oled_data = 16'b1100111011111110;
    else if (pixel_index == 3148 || pixel_index == 3340 || pixel_index == 3433) oled_data = 16'b1100011010111101;
    else if (pixel_index == 3149) oled_data = 16'b1011010111111010;
    else if (pixel_index == 3150) oled_data = 16'b1010010001001110;
    else if (pixel_index == 3151) oled_data = 16'b1001110100101100;
    else if (pixel_index == 3156) oled_data = 16'b0110001111001100;
    else if (pixel_index == 3162) oled_data = 16'b1000110110110110;
    else if (pixel_index == 3163 || pixel_index == 3638 || pixel_index == 4433 || pixel_index == 4436 || pixel_index == 4440 || pixel_index == 4581 || pixel_index == 4606) oled_data = 16'b1001011001111100;
    else if (pixel_index == 3165 || pixel_index == 3198 || pixel_index == 3235 || pixel_index == 3367 || pixel_index == 3546 || ((pixel_index >= 3574) && (pixel_index <= 3575)) || pixel_index == 3588 || ((pixel_index >= 3640) && (pixel_index <= 3647)) || pixel_index == 3742) oled_data = 16'b1001111001111101;
    else if (((pixel_index >= 3166) && (pixel_index <= 3167)) || pixel_index == 3631) oled_data = 16'b1001011000111101;
    else if (pixel_index == 3168) oled_data = 16'b0110110010111001;
    else if (pixel_index == 3170) oled_data = 16'b0101110011110111;
    else if (pixel_index == 3171) oled_data = 16'b0011001101001101;
    else if (pixel_index == 3174 || pixel_index == 5151) oled_data = 16'b1001110101110101;
    else if (pixel_index == 3175) oled_data = 16'b1010010111111000;
    else if (pixel_index == 3176 || pixel_index == 3248) oled_data = 16'b1000110000001011;
    else if (pixel_index == 3177) oled_data = 16'b1010010001001001;
    else if (pixel_index == 3178) oled_data = 16'b1010110011101011;
    else if (pixel_index == 3180) oled_data = 16'b1011010111110000;
    else if (pixel_index == 3181) oled_data = 16'b1011011001101110;
    else if (pixel_index == 3182) oled_data = 16'b1010111001101010;
    else if (pixel_index == 3183) oled_data = 16'b1011011000101101;
    else if (pixel_index == 3184) oled_data = 16'b1010011000101111;
    else if (pixel_index == 3185) oled_data = 16'b1010110111101100;
    else if (pixel_index == 3186 || pixel_index == 3188) oled_data = 16'b1011010111101001;
    else if (pixel_index == 3187) oled_data = 16'b1011011000100111;
    else if (pixel_index == 3190) oled_data = 16'b1000101111000101;
    else if (pixel_index == 3191) oled_data = 16'b1001110100110001;
    else if (pixel_index == 3192 || pixel_index == 4427) oled_data = 16'b1001010111111000;
    else if (pixel_index == 3193) oled_data = 16'b1010010111111010;
    else if (pixel_index == 3194 || pixel_index == 3328 || pixel_index == 3466 || pixel_index == 3672) oled_data = 16'b1010111001111011;
    else if (pixel_index == 3195) oled_data = 16'b1011111001111101;
    else if (pixel_index == 3196 || pixel_index == 3212 || pixel_index == 3384 || pixel_index == 3389 || pixel_index == 3487) oled_data = 16'b1011011010111110;
    else if (pixel_index == 3197 || pixel_index == 3454 || ((pixel_index >= 3481) && (pixel_index <= 3482)) || pixel_index == 3488 || ((pixel_index >= 3499) && (pixel_index <= 3500)) || ((pixel_index >= 3524) && (pixel_index <= 3525)) || ((pixel_index >= 3527) && (pixel_index <= 3528)) || pixel_index == 3583 || pixel_index == 3585 || pixel_index == 3690 || pixel_index == 4586) oled_data = 16'b1010111010111101;
    else if (pixel_index == 3199 || pixel_index == 3567 || pixel_index == 3590 || pixel_index == 3623 || ((pixel_index >= 3627) && (pixel_index <= 3628)) || pixel_index == 3675 || pixel_index == 3677 || pixel_index == 3717 || pixel_index == 3719 || pixel_index == 4567) oled_data = 16'b1010011001111101;
    else if (pixel_index == 3200) oled_data = 16'b1000110101110000;
    else if (pixel_index == 3201) oled_data = 16'b1001110101110010;
    else if (pixel_index == 3202 || pixel_index == 4439 || pixel_index == 4579) oled_data = 16'b1001111010111011;
    else if (pixel_index == 3203) oled_data = 16'b1001111100111101;
    else if (pixel_index == 3204 || pixel_index == 3632) oled_data = 16'b1000111010111101;
    else if (pixel_index == 3205) oled_data = 16'b1000011000111110;
    else if (pixel_index == 3206) oled_data = 16'b1000111000111110;
    else if (pixel_index == 3207 || pixel_index == 3660 || pixel_index == 3743) oled_data = 16'b1001111000111110;
    else if (pixel_index == 3208 || pixel_index == 3316 || pixel_index == 3383 || pixel_index == 3387 || pixel_index == 3396 || pixel_index == 3400 || pixel_index == 3438 || pixel_index == 3681 || pixel_index == 4573) oled_data = 16'b1011011010111101;
    else if (pixel_index == 3209) oled_data = 16'b1100011101111100;
    else if (pixel_index == 3210 || pixel_index == 3428) oled_data = 16'b1100011100111101;
    else if (pixel_index == 3211) oled_data = 16'b1011011011111110;
    else if (pixel_index == 3213) oled_data = 16'b1011111001111100;
    else if (pixel_index == 3214) oled_data = 16'b1101011101111110;
    else if (pixel_index == 3215) oled_data = 16'b0110101100001010;
    else if (pixel_index == 3216) oled_data = 16'b0010100011000011;
    else if (pixel_index == 3217) oled_data = 16'b0010100101000110;
    else if (pixel_index == 3218) oled_data = 16'b1001110111111011;
    else if (pixel_index == 3224) oled_data = 16'b0100101010001000;
    else if (pixel_index == 3231) oled_data = 16'b1010111000110111;
    else if (pixel_index == 3232 || pixel_index == 3602) oled_data = 16'b1011011011111111;
    else if (pixel_index == 3233 || pixel_index == 3450 || pixel_index == 3452 || pixel_index == 3483 || pixel_index == 3485 || pixel_index == 3617 || pixel_index == 4576) oled_data = 16'b1010111011111101;
    else if (pixel_index == 3236) oled_data = 16'b1011011001111101;
    else if (pixel_index == 3237 || pixel_index == 3295 || pixel_index == 4545) oled_data = 16'b1100111010111100;
    else if (pixel_index == 3238 || pixel_index == 3240 || pixel_index == 3259 || pixel_index == 3315 || pixel_index == 3334 || pixel_index == 4546 || pixel_index == 4549 || pixel_index == 4676 || pixel_index == 4678 || pixel_index == 4698 || pixel_index == 4877 || pixel_index == 5034) oled_data = 16'b1100111011111100;
    else if (pixel_index == 3239 || pixel_index == 4550 || pixel_index == 4685 || pixel_index == 4693 || pixel_index == 4700 || ((pixel_index >= 4702) && (pixel_index <= 4703)) || pixel_index == 5139 || pixel_index == 5710) oled_data = 16'b1100011010111011;
    else if (pixel_index == 3241 || pixel_index == 4695) oled_data = 16'b1100011011111100;
    else if (pixel_index == 3242 || pixel_index == 3329 || pixel_index == 3404 || pixel_index == 3453 || pixel_index == 3698 || pixel_index == 4553) oled_data = 16'b1011011010111100;
    else if (pixel_index == 3245) oled_data = 16'b1011111010111100;
    else if (pixel_index == 3246) oled_data = 16'b1010010110110101;
    else if (pixel_index == 3247 || pixel_index == 5516) oled_data = 16'b1010010100110011;
    else if (pixel_index == 3249) oled_data = 16'b1001010010101110;
    else if ((pixel_index >= 3250) && (pixel_index <= 3251)) oled_data = 16'b1010010101110011;
    else if (pixel_index == 3254) oled_data = 16'b1001010100101110;
    else if (pixel_index == 3256) oled_data = 16'b1011010110110000;
    else if (pixel_index == 3257 || pixel_index == 3285) oled_data = 16'b1011010111110011;
    else if (pixel_index == 3258 || pixel_index == 4538 || pixel_index == 5089 || pixel_index == 5129) oled_data = 16'b1011010111110111;
    else if (pixel_index == 3260) oled_data = 16'b1100111010111101;
    else if (pixel_index == 3261 || pixel_index == 3291 || pixel_index == 3336 || pixel_index == 3356 || pixel_index == 3391 || pixel_index == 3429 || pixel_index == 4547 || pixel_index == 4694 || pixel_index == 4697) oled_data = 16'b1100111011111101;
    else if (pixel_index == 3263 || pixel_index == 3301 || pixel_index == 3339 || pixel_index == 3341 || pixel_index == 3358 || pixel_index == 3430) oled_data = 16'b1011111011111101;
    else if (pixel_index == 3264) oled_data = 16'b0100101100001001;
    else if (pixel_index == 3265) oled_data = 16'b0011001000000110;
    else if (pixel_index == 3266) oled_data = 16'b0011001001001010;
    else if (pixel_index == 3271) oled_data = 16'b1000110110111001;
    else if (pixel_index == 3274) oled_data = 16'b1010110011101100;
    else if (pixel_index == 3275) oled_data = 16'b1011010100101100;
    else if (pixel_index == 3276) oled_data = 16'b1011010101101001;
    else if (pixel_index == 3277) oled_data = 16'b1011110111101000;
    else if (pixel_index == 3278) oled_data = 16'b1011010111100111;
    else if (pixel_index == 3279) oled_data = 16'b1011111001110000;
    else if (pixel_index == 3280) oled_data = 16'b1010111001110001;
    else if (pixel_index == 3282) oled_data = 16'b1011011000101110;
    else if (pixel_index == 3283) oled_data = 16'b1011110111101101;
    else if (pixel_index == 3284 || pixel_index == 3371) oled_data = 16'b1011110111110000;
    else if (pixel_index == 3286) oled_data = 16'b1010010100110000;
    else if (pixel_index == 3287 || pixel_index == 5334) oled_data = 16'b1010110111110111;
    else if (pixel_index == 3288 || pixel_index == 3354 || pixel_index == 3403 || pixel_index == 4692) oled_data = 16'b1011111010111011;
    else if (pixel_index == 3289 || pixel_index == 3292 || pixel_index == 3432) oled_data = 16'b1100011011111110;
    else if (pixel_index == 3293) oled_data = 16'b1100011010111110;
    else if (pixel_index == 3294 || pixel_index == 3394 || pixel_index == 3401) oled_data = 16'b1011111010111110;
    else if (pixel_index == 3296) oled_data = 16'b1011111000110011;
    else if (pixel_index == 3297 || (pixel_index >= 5348) && (pixel_index <= 5349)) oled_data = 16'b1100011010111001;
    else if (pixel_index == 3298 || pixel_index == 3300) oled_data = 16'b1100111100111110;
    else if (pixel_index == 3299 || pixel_index == 3303) oled_data = 16'b1100111101111110;
    else if (pixel_index == 3302) oled_data = 16'b1100111100111101;
    else if (pixel_index == 3304) oled_data = 16'b1101011011111110;
    else if (((pixel_index >= 3305) && (pixel_index <= 3306)) || pixel_index == 4661 || pixel_index == 4669 || pixel_index == 5492 || pixel_index == 5591) oled_data = 16'b1110011100111110;
    else if (pixel_index == 3307) oled_data = 16'b1101111100111110;
    else if (pixel_index == 3309 || (pixel_index >= 5010) && (pixel_index <= 5011)) oled_data = 16'b1101111101111100;
    else if (pixel_index == 3310 || pixel_index == 4541) oled_data = 16'b1100011001111001;
    else if (pixel_index == 3311 || pixel_index == 5327) oled_data = 16'b0100001000001000;
    else if (pixel_index == 3312) oled_data = 16'b0001100010000100;
    else if (pixel_index == 3313 || pixel_index == 4366) oled_data = 16'b0100101000001010;
    else if (pixel_index == 3314) oled_data = 16'b1101011101111101;
    else if (pixel_index == 3317) oled_data = 16'b1010110111111100;
    else if (pixel_index == 3318 || pixel_index == 3541 || pixel_index == 3598 || (pixel_index >= 4423) && (pixel_index <= 4424)) oled_data = 16'b1001010110111000;
    else if (pixel_index == 3322) oled_data = 16'b0011001000000001;
    else if (pixel_index == 3326) oled_data = 16'b0101101100000011;
    else if (pixel_index == 3327) oled_data = 16'b0111010000001100;
    else if (pixel_index == 3330 || pixel_index == 3414 || pixel_index == 3427 || pixel_index == 3451) oled_data = 16'b1011011011111101;
    else if (pixel_index == 3331 || pixel_index == 3386 || pixel_index == 3388 || pixel_index == 3390 || pixel_index == 3395 || pixel_index == 3434) oled_data = 16'b1011111011111110;
    else if (pixel_index == 3333 || pixel_index == 4666 || pixel_index == 4682) oled_data = 16'b1101011011111101;
    else if (pixel_index == 3337) oled_data = 16'b1100111010111110;
    else if (pixel_index == 3342 || pixel_index == 4555 || (pixel_index >= 4562) && (pixel_index <= 4563)) oled_data = 16'b1011011010111011;
    else if (pixel_index == 3343) oled_data = 16'b1010111001111000;
    else if (pixel_index == 3344) oled_data = 16'b1010110101110001;
    else if (pixel_index == 3345 || pixel_index == 5418 || pixel_index == 5880) oled_data = 16'b1011010110110100;
    else if (pixel_index == 3346 || pixel_index == 5056 || pixel_index == 5514) oled_data = 16'b1011110110110110;
    else if (pixel_index == 3347) oled_data = 16'b1100010111110100;
    else if ((pixel_index >= 3348) && (pixel_index <= 3349)) oled_data = 16'b1010110101110000;
    else if (pixel_index == 3350) oled_data = 16'b1010010110110010;
    else if (pixel_index == 3351) oled_data = 16'b1010110111110100;
    else if (pixel_index == 3352 || pixel_index == 3379) oled_data = 16'b1011111001110110;
    else if (pixel_index == 3353 || pixel_index == 3392 || pixel_index == 5363) oled_data = 16'b1011111001111010;
    else if (pixel_index == 3361 || pixel_index == 3746) oled_data = 16'b0100101010000110;
    else if (pixel_index == 3362) oled_data = 16'b0100001001001001;
    else if (pixel_index == 3363) oled_data = 16'b0110001111010000;
    else if (pixel_index == 3364 || pixel_index == 4613) oled_data = 16'b0110001111010001;
    else if (pixel_index == 3366) oled_data = 16'b1000010110110101;
    else if (pixel_index == 3368) oled_data = 16'b1000010111111000;
    else if (pixel_index == 3369) oled_data = 16'b1000110010110000;
    else if (pixel_index == 3370) oled_data = 16'b1011010110110011;
    else if (pixel_index == 3372) oled_data = 16'b1011010110101011;
    else if (pixel_index == 3373) oled_data = 16'b1011110111101100;
    else if (pixel_index == 3374) oled_data = 16'b1011111000101110;
    else if (pixel_index == 3375) oled_data = 16'b1011111001110100;
    else if (pixel_index == 3376) oled_data = 16'b1011111001110111;
    else if (((pixel_index >= 3377) && (pixel_index <= 3378)) || pixel_index == 3468) oled_data = 16'b1011011001110101;
    else if (pixel_index == 3380 || (pixel_index >= 5863) && (pixel_index <= 5864)) oled_data = 16'b1011011000110111;
    else if ((pixel_index >= 3381) && (pixel_index <= 3382)) oled_data = 16'b1010111001111010;
    else if (pixel_index == 3385 || pixel_index == 4561) oled_data = 16'b1011111100111110;
    else if (pixel_index == 3397) oled_data = 16'b1011111011111100;
    else if (pixel_index == 3398) oled_data = 16'b1011111100111100;
    else if (pixel_index == 3399) oled_data = 16'b1011011100111100;
    else if (pixel_index == 3405) oled_data = 16'b1100011101111110;
    else if (pixel_index == 3406 || pixel_index == 5351 || pixel_index == 6122) oled_data = 16'b1011110111111010;
    else if (pixel_index == 3407 || pixel_index == 5893 || pixel_index == 6057) oled_data = 16'b0110001101001110;
    else if (pixel_index == 3408 || pixel_index == 4559) oled_data = 16'b0011100110000110;
    else if (pixel_index == 3409) oled_data = 16'b0110101100001100;
    else if (pixel_index == 3410) oled_data = 16'b1011111100111101;
    else if (pixel_index == 3411) oled_data = 16'b1100011100111100;
    else if (pixel_index == 3413) oled_data = 16'b1100011011111111;
    else if (pixel_index == 3415) oled_data = 16'b1010011000111010;
    else if (pixel_index == 3416 || pixel_index == 5278) oled_data = 16'b1001010011110101;
    else if (pixel_index == 3417) oled_data = 16'b0110101111001110;
    else if (pixel_index == 3418) oled_data = 16'b0011101001000011;
    else if (pixel_index == 3423) oled_data = 16'b0111001110001001;
    else if (pixel_index == 3424) oled_data = 16'b1010010111110110;
    else if (pixel_index == 3425 || pixel_index == 3498) oled_data = 16'b1011011001111100;
    else if (pixel_index == 3440) oled_data = 16'b1010011000111000;
    else if ((pixel_index >= 3441) && (pixel_index <= 3442)) oled_data = 16'b1010111001111001;
    else if (pixel_index == 3443) oled_data = 16'b1011011000110110;
    else if (pixel_index == 3444 || pixel_index == 5858) oled_data = 16'b1010110110110101;
    else if (pixel_index == 3445) oled_data = 16'b1010010101110101;
    else if (pixel_index == 3446) oled_data = 16'b1010010110110110;
    else if (pixel_index == 3447 || pixel_index == 3539) oled_data = 16'b1010111000111000;
    else if (pixel_index == 3448 || (pixel_index >= 3471) && (pixel_index <= 3473)) oled_data = 16'b1010111000111010;
    else if (pixel_index == 3456) oled_data = 16'b0101001011000100;
    else if (pixel_index == 3458) oled_data = 16'b0100001000000011;
    else if (pixel_index == 3460) oled_data = 16'b0110001110001101;
    else if (pixel_index == 3463) oled_data = 16'b1000110111111000;
    else if (pixel_index == 3464) oled_data = 16'b1000010111111001;
    else if (pixel_index == 3465 || pixel_index == 3710) oled_data = 16'b1000110110110111;
    else if (pixel_index == 3467) oled_data = 16'b1011011010111000;
    else if (pixel_index == 3469) oled_data = 16'b1011011001110110;
    else if (pixel_index == 3470) oled_data = 16'b1011011010110111;
    else if (pixel_index == 3474) oled_data = 16'b1010011001111010;
    else if (pixel_index == 3475 || pixel_index == 4571) oled_data = 16'b1010011001111011;
    else if (pixel_index == 3476 || pixel_index == 4592) oled_data = 16'b1010011010111011;
    else if (((pixel_index >= 3478) && (pixel_index <= 3480)) || ((pixel_index >= 3521) && (pixel_index <= 3522)) || pixel_index == 3530 || pixel_index == 3547 || pixel_index == 3550 || pixel_index == 3564 || pixel_index == 3566 || ((pixel_index >= 3576) && (pixel_index <= 3577)) || pixel_index == 3580 || pixel_index == 3582 || pixel_index == 3604 || pixel_index == 3618 || pixel_index == 3622 || pixel_index == 3624 || pixel_index == 3629 || pixel_index == 3682 || pixel_index == 3689 || pixel_index == 3713 || ((pixel_index >= 3720) && (pixel_index <= 3721)) || pixel_index == 4583) oled_data = 16'b1010011010111101;
    else if (pixel_index == 3484 || pixel_index == 3494 || pixel_index == 3496 || pixel_index == 3531 || pixel_index == 3592 || pixel_index == 3716 || pixel_index == 4564 || pixel_index == 4577 || pixel_index == 4585 || (pixel_index >= 4599) && (pixel_index <= 4600)) oled_data = 16'b1010011010111100;
    else if (pixel_index == 3486 || pixel_index == 3506 || pixel_index == 3608) oled_data = 16'b1010111011111110;
    else if (pixel_index == 3489) oled_data = 16'b1010111010111111;
    else if (pixel_index == 3490 || pixel_index == 3508 || pixel_index == 3511 || pixel_index == 3526 || pixel_index == 3607 || pixel_index == 3621 || pixel_index == 3687) oled_data = 16'b1010111010111110;
    else if (pixel_index == 3491) oled_data = 16'b1001111000111100;
    else if (pixel_index == 3492 || pixel_index == 4565) oled_data = 16'b1010011000111100;
    else if (pixel_index == 3493 || pixel_index == 3537 || pixel_index == 3581 || pixel_index == 3684 || pixel_index == 3732 || pixel_index == 4575) oled_data = 16'b1010011011111101;
    else if (pixel_index == 3501) oled_data = 16'b1010111011111111;
    else if (pixel_index == 3502) oled_data = 16'b1001111000111010;
    else if (pixel_index == 3503) oled_data = 16'b0101101011001100;
    else if (pixel_index == 3504) oled_data = 16'b0011100101000100;
    else if (pixel_index == 3510 || pixel_index == 3630 || pixel_index == 3676 || pixel_index == 3718 || pixel_index == 3726 || pixel_index == 3741) oled_data = 16'b1001111001111110;
    else if (pixel_index == 3512 || pixel_index == 3659) oled_data = 16'b1001111000111101;
    else if (pixel_index == 3513) oled_data = 16'b0111110010110100;
    else if (pixel_index == 3514) oled_data = 16'b0100101001000011;
    else if (pixel_index == 3516) oled_data = 16'b0110110000001111;
    else if (pixel_index == 3520) oled_data = 16'b1001110110110101;
    else if (pixel_index == 3529 || pixel_index == 3532 || ((pixel_index >= 3699) && (pixel_index <= 3700)) || pixel_index == 3703 || pixel_index == 4572) oled_data = 16'b1010111001111100;
    else if (pixel_index == 3535 || pixel_index == 3544 || pixel_index == 3563 || pixel_index == 3587 || ((pixel_index >= 3625) && (pixel_index <= 3626)) || pixel_index == 3634 || ((pixel_index >= 4587) && (pixel_index <= 4588)) || pixel_index == 4593) oled_data = 16'b1001111001111100;
    else if (pixel_index == 3536 || pixel_index == 3639 || pixel_index == 3727 || pixel_index == 3736) oled_data = 16'b1001011010111101;
    else if (pixel_index == 3538) oled_data = 16'b1010011010111010;
    else if (pixel_index == 3540) oled_data = 16'b1001110110110111;
    else if (pixel_index == 3542 || ((pixel_index >= 4425) && (pixel_index <= 4426)) || pixel_index == 4429) oled_data = 16'b1001010111111001;
    else if (pixel_index == 3543 || ((pixel_index >= 4434) && (pixel_index <= 4435)) || pixel_index == 4438 || pixel_index == 4570) oled_data = 16'b1001011001111011;
    else if (pixel_index == 3552) oled_data = 16'b0101001011000010;
    else if (pixel_index == 3553) oled_data = 16'b0100101011000010;
    else if (pixel_index == 3562 || pixel_index == 3658 || pixel_index == 3731) oled_data = 16'b1001111001111011;
    else if (pixel_index == 3571 || pixel_index == 4590 || pixel_index == 4594 || pixel_index == 4597 || (pixel_index >= 4603) && (pixel_index <= 4604)) oled_data = 16'b1001111010111100;
    else if (pixel_index == 3579 || pixel_index == 3586 || pixel_index == 3701 || pixel_index == 4584) oled_data = 16'b1010011011111110;
    else if (pixel_index == 3589 || pixel_index == 4574) oled_data = 16'b1010011001111110;
    else if (pixel_index == 3591) oled_data = 16'b1010011000111101;
    else if (pixel_index == 3593 || pixel_index == 3664 || pixel_index == 4578) oled_data = 16'b1010011011111100;
    else if (pixel_index == 3595) oled_data = 16'b1010111001111110;
    else if (pixel_index == 3597 || pixel_index == 3723) oled_data = 16'b1010011010111111;
    else if (pixel_index == 3599 || pixel_index == 4271 || pixel_index == 4463) oled_data = 16'b0100000110000111;
    else if (pixel_index == 3601) oled_data = 16'b1000010110110111;
    else if (pixel_index == 3605 || pixel_index == 4437 || pixel_index == 4596) oled_data = 16'b1001011010111011;
    else if (pixel_index == 3606 || pixel_index == 3697) oled_data = 16'b1001111000111011;
    else if (pixel_index == 3609 || pixel_index == 4446 || pixel_index == 4448) oled_data = 16'b1000111000111010;
    else if (pixel_index == 3610) oled_data = 16'b0101101011000111;
    else if (pixel_index == 3611) oled_data = 16'b0110001100001010;
    else if (pixel_index == 3612 || pixel_index == 5794) oled_data = 16'b0111110001010000;
    else if (pixel_index == 3613 || pixel_index == 3615) oled_data = 16'b1000010011110001;
    else if (pixel_index == 3614) oled_data = 16'b0111110100110001;
    else if (pixel_index == 3616) oled_data = 16'b1001110111110110;
    else if (pixel_index == 3635) oled_data = 16'b1001111000111000;
    else if (((pixel_index >= 3636) && (pixel_index <= 3637)) || pixel_index == 4430) oled_data = 16'b1001011000111010;
    else if (pixel_index == 3648) oled_data = 16'b0110001100000000;
    else if (pixel_index == 3652) oled_data = 16'b0111110110110101;
    else if (pixel_index == 3656) oled_data = 16'b1000010001001110;
    else if (pixel_index == 3661) oled_data = 16'b1001111000111111;
    else if (pixel_index == 3663) oled_data = 16'b1001011011111110;
    else if ((pixel_index >= 3665) && (pixel_index <= 3666)) oled_data = 16'b1001111011111110;
    else if (pixel_index == 3670) oled_data = 16'b1010111001111111;
    else if (pixel_index == 3671) oled_data = 16'b1010111000111100;
    else if (pixel_index == 3673) oled_data = 16'b1010111000111101;
    else if (pixel_index == 3679 || pixel_index == 3704) oled_data = 16'b1010111011111011;
    else if (pixel_index == 3683 || pixel_index == 3686) oled_data = 16'b1010011011111111;
    else if (pixel_index == 3693 || pixel_index == 3734 || pixel_index == 4601) oled_data = 16'b1001111011111101;
    else if (pixel_index == 3694 || pixel_index == 4621) oled_data = 16'b0111010000010010;
    else if (pixel_index == 3695) oled_data = 16'b0011000011000100;
    else if (pixel_index == 3705 || ((pixel_index >= 4442) && (pixel_index <= 4443)) || pixel_index == 4607) oled_data = 16'b1000111001111100;
    else if (pixel_index == 3706 || pixel_index == 5135 || pixel_index == 5518) oled_data = 16'b0101101011001011;
    else if (pixel_index == 3709) oled_data = 16'b1001010011110010;
    else if (pixel_index == 3712) oled_data = 16'b1001111000110111;
    else if (pixel_index == 3724) oled_data = 16'b1001111001111111;
    else if (pixel_index == 3725) oled_data = 16'b1001011001111111;
    else if (pixel_index == 3728) oled_data = 16'b1000111011111110;
    else if (((pixel_index >= 3729) && (pixel_index <= 3730)) || pixel_index == 3740) oled_data = 16'b1001011001111101;
    else if (pixel_index == 3733) oled_data = 16'b1001011011111101;
    else if (pixel_index == 3744) oled_data = 16'b0101001011000001;
    else if (pixel_index == 3745) oled_data = 16'b0100101010000011;
    else if (pixel_index == 3749) oled_data = 16'b0101010100110110;
    else if (pixel_index == 3751) oled_data = 16'b0101110101111000;
    else if (pixel_index == 3752) oled_data = 16'b0101010110111010;
    else if (pixel_index == 3754 || pixel_index == 3765 || pixel_index == 3780 || pixel_index == 3794) oled_data = 16'b0110010111111100;
    else if (pixel_index == 3755 || pixel_index == 3785 || pixel_index == 3985) oled_data = 16'b0101110110111011;
    else if (pixel_index == 3756) oled_data = 16'b0110010110111001;
    else if (((pixel_index >= 3758) && (pixel_index <= 3762)) || pixel_index == 3773 || pixel_index == 3787 || pixel_index == 3798) oled_data = 16'b0110010111111011;
    else if (pixel_index == 3764) oled_data = 16'b0110010110111100;
    else if (pixel_index == 3766) oled_data = 16'b0110011001111101;
    else if (pixel_index == 3769 || pixel_index == 3772) oled_data = 16'b0110010111111010;
    else if (pixel_index == 3774 || pixel_index == 3783 || pixel_index == 4484 || pixel_index == 4487) oled_data = 16'b0110111000111011;
    else if (pixel_index == 3777 || pixel_index == 4182 || pixel_index == 4376 || pixel_index == 4454 || pixel_index == 4456) oled_data = 16'b0111011001111100;
    else if (pixel_index == 3786 || pixel_index == 3796 || pixel_index == 3828) oled_data = 16'b0101110110111010;
    else if (pixel_index == 3789 || pixel_index == 4323) oled_data = 16'b0101010101111000;
    else if (pixel_index == 3790 || pixel_index == 5981) oled_data = 16'b0011101001001010;
    else if (pixel_index == 3791) oled_data = 16'b0010000011000011;
    else if (pixel_index == 3793 || pixel_index == 3827) oled_data = 16'b0101110101111001;
    else if (pixel_index == 3800) oled_data = 16'b0110010011110111;
    else if (pixel_index == 3801 || pixel_index == 3804) oled_data = 16'b0101110001010000;
    else if (pixel_index == 3802) oled_data = 16'b0100101101001011;
    else if (pixel_index == 3803) oled_data = 16'b0101110000001111;
    else if (pixel_index == 3805) oled_data = 16'b0101101111001101;
    else if (pixel_index == 3807) oled_data = 16'b0101001111010011;
    else if (pixel_index == 3808) oled_data = 16'b0101010010110110;
    else if (((pixel_index >= 3810) && (pixel_index <= 3811)) || pixel_index == 3815) oled_data = 16'b0101010011111001;
    else if (pixel_index == 3813) oled_data = 16'b0101110011111001;
    else if (pixel_index == 3818) oled_data = 16'b0101010100111001;
    else if (pixel_index == 3819 || pixel_index == 3834 || pixel_index == 3836 || (pixel_index >= 3838) && (pixel_index <= 3839)) oled_data = 16'b0101110101111010;
    else if (pixel_index == 3820 || pixel_index == 3829) oled_data = 16'b0101110100111001;
    else if (pixel_index == 3821) oled_data = 16'b0101010101111001;
    else if (pixel_index == 3822) oled_data = 16'b0101110110111001;
    else if (pixel_index == 3824) oled_data = 16'b0101010011111010;
    else if (pixel_index == 3826 || pixel_index == 3830 || pixel_index == 3837) oled_data = 16'b0101110100111010;
    else if (pixel_index == 3832) oled_data = 16'b0101110100111011;
    else if (pixel_index == 3833) oled_data = 16'b0101110011111010;
    else if (pixel_index == 3840) oled_data = 16'b0100101011000011;
    else if (pixel_index == 3842) oled_data = 16'b0010101001000111;
    else if (pixel_index == 3843) oled_data = 16'b0010001010001000;
    else if (pixel_index == 3845) oled_data = 16'b0001010000010101;
    else if (pixel_index == 3846) oled_data = 16'b0000110000011000;
    else if (pixel_index == 3847 || ((pixel_index >= 3855) && (pixel_index <= 3856)) || pixel_index == 3858 || ((pixel_index >= 3928) && (pixel_index <= 3929)) || pixel_index == 3942) oled_data = 16'b0000110010111000;
    else if (((pixel_index >= 3848) && (pixel_index <= 3849)) || pixel_index == 3940 || pixel_index == 3944 || pixel_index == 3949) oled_data = 16'b0001010010111001;
    else if (pixel_index == 3850 || pixel_index == 3854 || (pixel_index >= 3859) && (pixel_index <= 3860)) oled_data = 16'b0000110010111001;
    else if (pixel_index == 3851) oled_data = 16'b0000010010111000;
    else if (pixel_index == 3852) oled_data = 16'b0000110010110111;
    else if (pixel_index == 3853) oled_data = 16'b0000110001010111;
    else if (pixel_index == 3857 || pixel_index == 3923) oled_data = 16'b0001010010111000;
    else if (pixel_index == 3861 || pixel_index == 3866 || ((pixel_index >= 3930) && (pixel_index <= 3932)) || pixel_index == 3945 || pixel_index == 3950) oled_data = 16'b0001010011111000;
    else if ((pixel_index >= 3862) && (pixel_index <= 3863)) oled_data = 16'b0001010011111001;
    else if (pixel_index == 3864) oled_data = 16'b0001010011111010;
    else if (pixel_index == 3865 || pixel_index == 3951) oled_data = 16'b0001110011111001;
    else if (pixel_index == 3867) oled_data = 16'b0001110011111010;
    else if (pixel_index == 3868) oled_data = 16'b0001110100111000;
    else if (((pixel_index >= 3869) && (pixel_index <= 3870)) || pixel_index == 3959) oled_data = 16'b0010010100111001;
    else if (pixel_index == 3871) oled_data = 16'b0001110100111010;
    else if (pixel_index == 3872 || pixel_index == 3955 || pixel_index == 3958 || pixel_index == 4018) oled_data = 16'b0010010100111010;
    else if (pixel_index == 3873) oled_data = 16'b0010010101111010;
    else if (pixel_index == 3874) oled_data = 16'b0010010100110111;
    else if (pixel_index == 3875) oled_data = 16'b0010010011111000;
    else if (pixel_index == 3876) oled_data = 16'b0010010011111010;
    else if (((pixel_index >= 3877) && (pixel_index <= 3878)) || pixel_index == 4011) oled_data = 16'b0010010011111001;
    else if (pixel_index == 3880) oled_data = 16'b0011010100111000;
    else if (pixel_index == 3881 || pixel_index == 3892 || pixel_index == 3970) oled_data = 16'b0011010100111001;
    else if (pixel_index == 3882 || pixel_index == 3894 || pixel_index == 3963 || (pixel_index >= 3965) && (pixel_index <= 3966)) oled_data = 16'b0011010101111010;
    else if ((pixel_index >= 3883) && (pixel_index <= 3884)) oled_data = 16'b0011110110111011;
    else if (pixel_index == 3885) oled_data = 16'b0100110000010101;
    else if (pixel_index == 3886) oled_data = 16'b0011101000001000;
    else if (pixel_index == 3888 || pixel_index == 4513) oled_data = 16'b0010000110000111;
    else if (pixel_index == 3889 || pixel_index == 3971) oled_data = 16'b0011110100111010;
    else if (pixel_index == 3890) oled_data = 16'b0011110101111010;
    else if (pixel_index == 3900) oled_data = 16'b0011101111001111;
    else if (pixel_index == 3901) oled_data = 16'b0100001110001100;
    else if (pixel_index == 3904) oled_data = 16'b0011110001010111;
    else if (pixel_index == 3907) oled_data = 16'b0011001111011000;
    else if (((pixel_index >= 3908) && (pixel_index <= 3909)) || pixel_index == 4006 || pixel_index == 4008) oled_data = 16'b0010010000010111;
    else if (pixel_index == 3910) oled_data = 16'b0001110000010111;
    else if (pixel_index == 3914) oled_data = 16'b0001110000010110;
    else if (pixel_index == 3915) oled_data = 16'b0001110001011000;
    else if (pixel_index == 3916 || pixel_index == 3922 || pixel_index == 3925 || pixel_index == 3943) oled_data = 16'b0001010010110111;
    else if (pixel_index == 3917) oled_data = 16'b0001110010110111;
    else if (pixel_index == 3918) oled_data = 16'b0001010011110111;
    else if (pixel_index == 3919 || pixel_index == 3921 || pixel_index == 3927) oled_data = 16'b0001010001011000;
    else if (pixel_index == 3924 || (pixel_index >= 4013) && (pixel_index <= 4014)) oled_data = 16'b0001110011111000;
    else if (pixel_index == 3926) oled_data = 16'b0001010001010111;
    else if (pixel_index == 3933 || pixel_index == 3935 || pixel_index == 3953) oled_data = 16'b0001010100111001;
    else if (pixel_index == 3934) oled_data = 16'b0000110100111001;
    else if (pixel_index == 3937) oled_data = 16'b0011001101001011;
    else if (pixel_index == 3938) oled_data = 16'b0010001111010001;
    else if (pixel_index == 3939) oled_data = 16'b0001110000010100;
    else if (pixel_index == 3941) oled_data = 16'b0000110010111010;
    else if (pixel_index == 3946) oled_data = 16'b0000110011111001;
    else if (pixel_index == 3947) oled_data = 16'b0000110011111010;
    else if (pixel_index == 3948) oled_data = 16'b0000010011111000;
    else if (pixel_index == 3952) oled_data = 16'b0001010100111000;
    else if (pixel_index == 3954 || ((pixel_index >= 4021) && (pixel_index <= 4025)) || pixel_index == 4035) oled_data = 16'b0001110101111000;
    else if (pixel_index == 3956) oled_data = 16'b0001110100111001;
    else if (pixel_index == 3960 || pixel_index == 3962 || pixel_index == 3967) oled_data = 16'b0010110100111001;
    else if (pixel_index == 3961 || pixel_index == 3964) oled_data = 16'b0011010100111010;
    else if ((pixel_index >= 3968) && (pixel_index <= 3969)) oled_data = 16'b0010110101111010;
    else if (pixel_index == 3972) oled_data = 16'b0100010101111010;
    else if (pixel_index == 3973 || pixel_index == 4059) oled_data = 16'b0100010110111010;
    else if (pixel_index == 3974) oled_data = 16'b0100010101111001;
    else if (pixel_index == 3975) oled_data = 16'b0100110110111001;
    else if (pixel_index == 3976 || pixel_index == 3980) oled_data = 16'b0101010110111001;
    else if (pixel_index == 3977) oled_data = 16'b0100110110111010;
    else if (pixel_index == 3979) oled_data = 16'b0100110110111011;
    else if (pixel_index == 3981 || pixel_index == 4077) oled_data = 16'b0110010001010101;
    else if (pixel_index == 3982) oled_data = 16'b0100101000001001;
    else if (pixel_index == 3984 || pixel_index == 5985 || pixel_index == 5987) oled_data = 16'b0011001000001001;
    else if (pixel_index == 3988) oled_data = 16'b0110010100111001;
    else if (pixel_index == 3989) oled_data = 16'b0110010101111100;
    else if (pixel_index == 3990) oled_data = 16'b0101110111111010;
    else if (pixel_index == 3991) oled_data = 16'b0110010011110110;
    else if (pixel_index == 3994 || pixel_index == 4995 || pixel_index == 4997) oled_data = 16'b0110001101001111;
    else if (pixel_index == 3998) oled_data = 16'b0100010010110111;
    else if (pixel_index == 4005) oled_data = 16'b0011010001010111;
    else if (pixel_index == 4007) oled_data = 16'b0010010000011000;
    else if (pixel_index == 4010) oled_data = 16'b0010010010111001;
    else if (pixel_index == 4012) oled_data = 16'b0001110010111001;
    else if (pixel_index == 4015) oled_data = 16'b0010010010111000;
    else if (pixel_index == 4016) oled_data = 16'b0010110011111000;
    else if (pixel_index == 4017) oled_data = 16'b0010010100111000;
    else if (pixel_index == 4019) oled_data = 16'b0001110110111010;
    else if (pixel_index == 4020) oled_data = 16'b0010010101111001;
    else if (pixel_index == 4026) oled_data = 16'b0010010110111001;
    else if (pixel_index == 4027 || ((pixel_index >= 4049) && (pixel_index <= 4050)) || pixel_index == 4052) oled_data = 16'b0010010111111010;
    else if (pixel_index == 4028 || pixel_index == 4030 || pixel_index == 4048) oled_data = 16'b0001110110111001;
    else if (pixel_index == 4029 || pixel_index == 4031 || ((pixel_index >= 4039) && (pixel_index <= 4040)) || (pixel_index >= 4045) && (pixel_index <= 4047)) oled_data = 16'b0001110111111010;
    else if (pixel_index == 4032) oled_data = 16'b0100110000001011;
    else if (pixel_index == 4033) oled_data = 16'b0011110010110000;
    else if (pixel_index == 4034) oled_data = 16'b0010110011110101;
    else if (pixel_index == 4036) oled_data = 16'b0001010110111011;
    else if (pixel_index == 4037) oled_data = 16'b0001010111111100;
    else if (pixel_index == 4038) oled_data = 16'b0001011000111010;
    else if (pixel_index == 4041) oled_data = 16'b0001110111111001;
    else if (pixel_index == 4042) oled_data = 16'b0000111000111010;
    else if (pixel_index == 4043) oled_data = 16'b0000110111111010;
    else if (pixel_index == 4044) oled_data = 16'b0001010110111001;
    else if (pixel_index == 4051 || ((pixel_index >= 4054) && (pixel_index <= 4055)) || pixel_index == 4132) oled_data = 16'b0010110111111010;
    else if (pixel_index == 4053) oled_data = 16'b0010110101111001;
    else if (pixel_index == 4056) oled_data = 16'b0011010111111010;
    else if (pixel_index == 4057) oled_data = 16'b0011010111111011;
    else if (pixel_index == 4058 || pixel_index == 4063 || pixel_index == 4065) oled_data = 16'b0011110110111010;
    else if (pixel_index == 4060 || pixel_index == 4062 || pixel_index == 4327) oled_data = 16'b0100010111111011;
    else if (pixel_index == 4061) oled_data = 16'b0100010110111100;
    else if (pixel_index == 4064) oled_data = 16'b0011110111111011;
    else if (pixel_index == 4066) oled_data = 16'b0100010101111011;
    else if (pixel_index == 4067) oled_data = 16'b0100010111111100;
    else if (pixel_index == 4068 || pixel_index == 4103 || pixel_index == 4156 || pixel_index == 4331 || (pixel_index >= 4337) && (pixel_index <= 4338)) oled_data = 16'b0100011000111011;
    else if (pixel_index == 4069 || pixel_index == 4101) oled_data = 16'b0100011001111010;
    else if (pixel_index == 4070 || pixel_index == 4099 || pixel_index == 4155 || pixel_index == 4341 || pixel_index == 4347 || (pixel_index >= 4349) && (pixel_index <= 4350)) oled_data = 16'b0100111000111011;
    else if (pixel_index == 4071 || pixel_index == 4343 || pixel_index == 4391) oled_data = 16'b0101011000111011;
    else if (((pixel_index >= 4072) && (pixel_index <= 4073)) || pixel_index == 4097 || pixel_index == 4161 || pixel_index == 4261 || pixel_index == 4286 || pixel_index == 4291 || pixel_index == 4345 || pixel_index == 4480) oled_data = 16'b0101111001111100;
    else if (pixel_index == 4074 || pixel_index == 4157 || pixel_index == 4392) oled_data = 16'b0101011000111100;
    else if (pixel_index == 4075) oled_data = 16'b0101111000111100;
    else if (pixel_index == 4076 || pixel_index == 4098 || pixel_index == 4389) oled_data = 16'b0101011001111011;
    else if (pixel_index == 4078 || pixel_index == 4270) oled_data = 16'b0110001010001011;
    else if (pixel_index == 4081 || pixel_index == 4086 || pixel_index == 4167 || pixel_index == 4169 || pixel_index == 4257 || pixel_index == 4260 || pixel_index == 4288 || pixel_index == 4385 || pixel_index == 4497 || pixel_index == 4499 || pixel_index == 4506 || pixel_index == 4509) oled_data = 16'b0110011010111100;
    else if (pixel_index == 4082 || pixel_index == 4096 || pixel_index == 4466) oled_data = 16'b0110011001111100;
    else if (pixel_index == 4083 || pixel_index == 4355) oled_data = 16'b0101111010111011;
    else if (pixel_index == 4084) oled_data = 16'b0101111000111011;
    else if (pixel_index == 4085 || pixel_index == 4171 || pixel_index == 4181 || pixel_index == 4195 || pixel_index == 4501) oled_data = 16'b0101111010111101;
    else if (pixel_index == 4087) oled_data = 16'b0110110111111000;
    else if (pixel_index == 4088) oled_data = 16'b0110110101110101;
    else if (pixel_index == 4090) oled_data = 16'b0110110100110100;
    else if (pixel_index == 4091) oled_data = 16'b0101110110110100;
    else if (pixel_index == 4093) oled_data = 16'b0101110101110100;
    else if (pixel_index == 4094) oled_data = 16'b0101111000111010;
    else if (pixel_index == 4095 || pixel_index == 4386) oled_data = 16'b0110111010111011;
    else if (pixel_index == 4100) oled_data = 16'b0100011000111010;
    else if (pixel_index == 4102 || pixel_index == 4145 || pixel_index == 4242 || pixel_index == 4247 || pixel_index == 4250 || pixel_index == 4295) oled_data = 16'b0011111001111011;
    else if (pixel_index == 4104 || pixel_index == 4333) oled_data = 16'b0011111000111100;
    else if (pixel_index == 4105 || pixel_index == 4208 || pixel_index == 4303) oled_data = 16'b0011011010111100;
    else if (pixel_index == 4106 || pixel_index == 4294 || pixel_index == 4310 || ((pixel_index >= 4316) && (pixel_index <= 4317)) || ((pixel_index >= 4329) && (pixel_index <= 4330)) || pixel_index == 4399) oled_data = 16'b0011111001111100;
    else if (pixel_index == 4107 || pixel_index == 4240) oled_data = 16'b0011011011111100;
    else if (pixel_index == 4108 || pixel_index == 4233) oled_data = 16'b0010111010111100;
    else if (pixel_index == 4109 || pixel_index == 4211 || pixel_index == 4219 || pixel_index == 4234 || pixel_index == 4402) oled_data = 16'b0010011010111100;
    else if (pixel_index == 4110 || ((pixel_index >= 4118) && (pixel_index <= 4120)) || pixel_index == 4213 || pixel_index == 4235) oled_data = 16'b0001111010111011;
    else if (pixel_index == 4111 || pixel_index == 4141 || pixel_index == 4144 || pixel_index == 4153) oled_data = 16'b0011011000111010;
    else if (pixel_index == 4112 || pixel_index == 4245 || (pixel_index >= 4335) && (pixel_index <= 4336)) oled_data = 16'b0011011001111011;
    else if (pixel_index == 4113) oled_data = 16'b0010111010111011;
    else if (pixel_index == 4114 || pixel_index == 4122 || pixel_index == 4215 || (pixel_index >= 4217) && (pixel_index <= 4218)) oled_data = 16'b0001111011111100;
    else if (pixel_index == 4115 || pixel_index == 4126) oled_data = 16'b0001011011111101;
    else if (pixel_index == 4116) oled_data = 16'b0001011010111101;
    else if (pixel_index == 4117 || pixel_index == 4124) oled_data = 16'b0001011011111100;
    else if (pixel_index == 4121) oled_data = 16'b0001111011111011;
    else if (pixel_index == 4123) oled_data = 16'b0010011011111100;
    else if (pixel_index == 4125) oled_data = 16'b0001111100111100;
    else if (pixel_index == 4127) oled_data = 16'b0001011100111101;
    else if (pixel_index == 4130) oled_data = 16'b0011110001010001;
    else if (pixel_index == 4131) oled_data = 16'b0010010101110101;
    else if (pixel_index == 4133 || pixel_index == 4136 || pixel_index == 4140 || pixel_index == 4147 || (pixel_index >= 4230) && (pixel_index <= 4231)) oled_data = 16'b0010011000111010;
    else if (pixel_index == 4134) oled_data = 16'b0010011000111001;
    else if (pixel_index == 4135) oled_data = 16'b0010010111111000;
    else if (pixel_index == 4137 || pixel_index == 4148) oled_data = 16'b0010111000111010;
    else if (pixel_index == 4138) oled_data = 16'b0010011001111011;
    else if (pixel_index == 4139) oled_data = 16'b0001111000111011;
    else if (pixel_index == 4142) oled_data = 16'b0011011001111001;
    else if (pixel_index == 4143 || pixel_index == 4152) oled_data = 16'b0011011001111010;
    else if (pixel_index == 4146) oled_data = 16'b0010111000111011;
    else if (pixel_index == 4149) oled_data = 16'b0010011000111011;
    else if (pixel_index == 4150 || pixel_index == 4232 || pixel_index == 4244 || ((pixel_index >= 4305) && (pixel_index <= 4306)) || pixel_index == 4312 || pixel_index == 4401) oled_data = 16'b0010111001111100;
    else if (pixel_index == 4151) oled_data = 16'b0010111001111011;
    else if (pixel_index == 4154 || pixel_index == 4334) oled_data = 16'b0011011000111011;
    else if (pixel_index == 4158 || pixel_index == 4170 || pixel_index == 4287 || pixel_index == 4346 || pixel_index == 4390) oled_data = 16'b0101011001111100;
    else if (pixel_index == 4159 || pixel_index == 4353) oled_data = 16'b0101011001111010;
    else if (pixel_index == 4160 || pixel_index == 4289 || pixel_index == 4384 || pixel_index == 4467 || pixel_index == 4479 || pixel_index == 4496) oled_data = 16'b0110011010111101;
    else if (((pixel_index >= 4162) && (pixel_index <= 4163)) || pixel_index == 4344) oled_data = 16'b0110011000111100;
    else if (pixel_index == 4164 || pixel_index == 4166 || pixel_index == 4255 || pixel_index == 4262 || pixel_index == 4267 || pixel_index == 4504 || pixel_index == 4508) oled_data = 16'b0101111010111100;
    else if (pixel_index == 4165 || pixel_index == 4179 || pixel_index == 4263) oled_data = 16'b0101011010111100;
    else if (pixel_index == 4168 || pixel_index == 4172 || pixel_index == 4268 || pixel_index == 4277 || pixel_index == 4491 || pixel_index == 4494) oled_data = 16'b0110111010111100;
    else if (pixel_index == 4173) oled_data = 16'b0111110100110111;
    else if (pixel_index == 4174) oled_data = 16'b0111101100001100;
    else if (pixel_index == 4175) oled_data = 16'b0101001001001000;
    else if (pixel_index == 4177) oled_data = 16'b0101111011111110;
    else if (pixel_index == 4178 || pixel_index == 4478 || pixel_index == 4485 || pixel_index == 4490 || pixel_index == 4492) oled_data = 16'b0110111001111100;
    else if (pixel_index == 4180 || pixel_index == 4388 || (pixel_index >= 4481) && (pixel_index <= 4482)) oled_data = 16'b0101111001111011;
    else if (pixel_index == 4183) oled_data = 16'b0111011000111010;
    else if (pixel_index == 4185) oled_data = 16'b0111110111111000;
    else if (pixel_index == 4186) oled_data = 16'b1000110101111000;
    else if (pixel_index == 4187) oled_data = 16'b0111011000111000;
    else if (pixel_index == 4188) oled_data = 16'b0110111000111000;
    else if (pixel_index == 4189) oled_data = 16'b0111111000110111;
    else if (pixel_index == 4190) oled_data = 16'b0111111011111100;
    else if (pixel_index == 4191) oled_data = 16'b1000011011111100;
    else if (pixel_index == 4192) oled_data = 16'b0111111011111101;
    else if (pixel_index == 4193 || pixel_index == 4371) oled_data = 16'b0111011011111101;
    else if (pixel_index == 4194 || pixel_index == 4256 || pixel_index == 4276 || pixel_index == 4498 || pixel_index == 4500) oled_data = 16'b0110011011111101;
    else if (pixel_index == 4196) oled_data = 16'b0101011011111101;
    else if (pixel_index == 4197) oled_data = 16'b0101011011111100;
    else if (pixel_index == 4198 || pixel_index == 4362 || pixel_index == 4507) oled_data = 16'b0101111011111100;
    else if ((pixel_index >= 4199) && (pixel_index <= 4200)) oled_data = 16'b0101111100111101;
    else if (pixel_index == 4201) oled_data = 16'b0100011011111101;
    else if ((pixel_index >= 4202) && (pixel_index <= 4203)) oled_data = 16'b0100111100111101;
    else if (pixel_index == 4204) oled_data = 16'b0100011100111101;
    else if (pixel_index == 4205 || pixel_index == 4293 || pixel_index == 4299 || pixel_index == 4308 || pixel_index == 4406) oled_data = 16'b0100011010111100;
    else if (pixel_index == 4206 || ((pixel_index >= 4248) && (pixel_index <= 4249)) || pixel_index == 4319 || pixel_index == 4360 || pixel_index == 4408) oled_data = 16'b0011111010111100;
    else if (pixel_index == 4207) oled_data = 16'b0011111011111100;
    else if ((pixel_index >= 4209) && (pixel_index <= 4210)) oled_data = 16'b0010111011111100;
    else if (pixel_index == 4212 || pixel_index == 4216 || (pixel_index >= 4220) && (pixel_index <= 4222)) oled_data = 16'b0001111010111100;
    else if (pixel_index == 4214) oled_data = 16'b0001011011111011;
    else if (pixel_index == 4223) oled_data = 16'b0001011010111100;
    else if (pixel_index == 4225) oled_data = 16'b0101110010101110;
    else if (pixel_index == 4226) oled_data = 16'b0100110001001111;
    else if (pixel_index == 4227) oled_data = 16'b0100110011110000;
    else if (pixel_index == 4228) oled_data = 16'b0100010101110100;
    else if (pixel_index == 4229) oled_data = 16'b0010110111110111;
    else if (pixel_index == 4236 || pixel_index == 4238) oled_data = 16'b0010011010111011;
    else if (pixel_index == 4237) oled_data = 16'b0010011010111010;
    else if (pixel_index == 4239) oled_data = 16'b0010111010111010;
    else if (pixel_index == 4241 || pixel_index == 4309) oled_data = 16'b0011111010111011;
    else if (pixel_index == 4243 || pixel_index == 4313 || pixel_index == 4332) oled_data = 16'b0011011000111100;
    else if (pixel_index == 4246 || pixel_index == 4307) oled_data = 16'b0011011010111011;
    else if (pixel_index == 4251 || ((pixel_index >= 4296) && (pixel_index <= 4298)) || ((pixel_index >= 4314) && (pixel_index <= 4315)) || pixel_index == 4318 || ((pixel_index >= 4396) && (pixel_index <= 4397)) || pixel_index == 4404 || pixel_index == 4407 || pixel_index == 4412) oled_data = 16'b0100011001111100;
    else if (pixel_index == 4252 || pixel_index == 4265 || pixel_index == 4300) oled_data = 16'b0100011010111011;
    else if (pixel_index == 4253) oled_data = 16'b0100011001111011;
    else if (pixel_index == 4254 || pixel_index == 4264 || pixel_index == 4409 || pixel_index == 4413) oled_data = 16'b0100111010111100;
    else if ((pixel_index >= 4258) && (pixel_index <= 4259)) oled_data = 16'b0110011010111011;
    else if (pixel_index == 4266 || pixel_index == 4356) oled_data = 16'b0101011010111011;
    else if (pixel_index == 4269 || pixel_index == 5064) oled_data = 16'b1000110100110011;
    else if (pixel_index == 4273) oled_data = 16'b0110111100111101;
    else if (pixel_index == 4274 || pixel_index == 4372) oled_data = 16'b0111011011111110;
    else if (pixel_index == 4275) oled_data = 16'b0110111011111110;
    else if (pixel_index == 4278) oled_data = 16'b1000111010111100;
    else if (pixel_index == 4279 || pixel_index == 4380 || pixel_index == 4457) oled_data = 16'b0111011010111101;
    else if (pixel_index == 4280 || pixel_index == 4468) oled_data = 16'b0111011001111101;
    else if (pixel_index == 4281 || pixel_index == 4364) oled_data = 16'b0111011001111010;
    else if (pixel_index == 4282) oled_data = 16'b0110111000111001;
    else if (pixel_index == 4283) oled_data = 16'b0110011001111010;
    else if (pixel_index == 4284) oled_data = 16'b0101111001111010;
    else if (pixel_index == 4285) oled_data = 16'b0101011000111001;
    else if (pixel_index == 4290 || pixel_index == 4410 || pixel_index == 4503) oled_data = 16'b0101011010111101;
    else if (pixel_index == 4292 || pixel_index == 4351 || pixel_index == 4359 || pixel_index == 4395 || pixel_index == 4411) oled_data = 16'b0100111001111100;
    else if (pixel_index == 4301) oled_data = 16'b0100111010111011;
    else if (pixel_index == 4302) oled_data = 16'b0100111011111011;
    else if (pixel_index == 4304) oled_data = 16'b0011011001111101;
    else if (pixel_index == 4311) oled_data = 16'b0011011001111100;
    else if (pixel_index == 4321) oled_data = 16'b0011110011110111;
    else if (pixel_index == 4322) oled_data = 16'b0011110101111000;
    else if (pixel_index == 4324) oled_data = 16'b0100110111111000;
    else if (pixel_index == 4325) oled_data = 16'b0011110111111010;
    else if (pixel_index == 4326 || (pixel_index >= 4339) && (pixel_index <= 4340)) oled_data = 16'b0011111000111011;
    else if (pixel_index == 4328) oled_data = 16'b0100111000111100;
    else if (pixel_index == 4342) oled_data = 16'b0101011000111010;
    else if (pixel_index == 4348 || pixel_index == 4352 || (pixel_index >= 4357) && (pixel_index <= 4358)) oled_data = 16'b0100111001111011;
    else if (pixel_index == 4354 || (pixel_index >= 4393) && (pixel_index <= 4394)) oled_data = 16'b0100111001111101;
    else if (pixel_index == 4361) oled_data = 16'b0100011010111101;
    else if (pixel_index == 4363 || pixel_index == 4379) oled_data = 16'b0111011011111100;
    else if (pixel_index == 4365 || pixel_index == 4531) oled_data = 16'b0111010001010001;
    else if (pixel_index == 4367) oled_data = 16'b0011000110000111;
    else if (pixel_index == 4369) oled_data = 16'b1000011101111100;
    else if (pixel_index == 4370 || pixel_index == 4510) oled_data = 16'b0110011011111100;
    else if (pixel_index == 4373) oled_data = 16'b1000011011111110;
    else if (pixel_index == 4374) oled_data = 16'b1001011011111100;
    else if (pixel_index == 4375) oled_data = 16'b1000011011111101;
    else if (pixel_index == 4377) oled_data = 16'b0111111001111011;
    else if (pixel_index == 4378) oled_data = 16'b0111111001111101;
    else if (pixel_index == 4381 || pixel_index == 4489) oled_data = 16'b0110111001111101;
    else if (pixel_index == 4382) oled_data = 16'b0110111010111110;
    else if (pixel_index == 4383) oled_data = 16'b0110011011111110;
    else if (pixel_index == 4387 || pixel_index == 4470 || pixel_index == 4486 || pixel_index == 4493) oled_data = 16'b0110111001111011;
    else if (pixel_index == 4398) oled_data = 16'b0100011000111100;
    else if (pixel_index == 4400) oled_data = 16'b0011111001111101;
    else if (pixel_index == 4403) oled_data = 16'b0011011010111101;
    else if (pixel_index == 4405) oled_data = 16'b0100111010111101;
    else if (pixel_index == 4414) oled_data = 16'b0101011001111101;
    else if (pixel_index == 4415) oled_data = 16'b0101111001111101;
    else if (pixel_index == 4416 || pixel_index == 4614) oled_data = 16'b0110110000010011;
    else if (pixel_index == 4419) oled_data = 16'b1000010011110110;
    else if (pixel_index == 4420) oled_data = 16'b1000110011110111;
    else if (pixel_index == 4421) oled_data = 16'b1000110101110111;
    else if (pixel_index == 4422) oled_data = 16'b1000110110111000;
    else if (pixel_index == 4428) oled_data = 16'b1001010111111010;
    else if ((pixel_index >= 4431) && (pixel_index <= 4432)) oled_data = 16'b1000111000111100;
    else if (pixel_index == 4441 || pixel_index == 4580 || pixel_index == 4595 || pixel_index == 4605) oled_data = 16'b1001011010111100;
    else if ((pixel_index >= 4444) && (pixel_index <= 4445)) oled_data = 16'b1000011000111011;
    else if (pixel_index == 4449) oled_data = 16'b1000010111111010;
    else if (pixel_index == 4451 || pixel_index == 4455 || pixel_index == 4474) oled_data = 16'b0111111001111100;
    else if ((pixel_index >= 4452) && (pixel_index <= 4453)) oled_data = 16'b0111111001111010;
    else if (pixel_index == 4458) oled_data = 16'b1000011001111011;
    else if (pixel_index == 4459) oled_data = 16'b1000011001111100;
    else if (pixel_index == 4461) oled_data = 16'b0110001111001111;
    else if (pixel_index == 4462 || (pixel_index >= 5888) && (pixel_index <= 5889)) oled_data = 16'b0100001000001001;
    else if (pixel_index == 4465) oled_data = 16'b0111011010111011;
    else if (pixel_index == 4469) oled_data = 16'b0111111010111011;
    else if (pixel_index == 4473) oled_data = 16'b0111011001111011;
    else if (pixel_index == 4475) oled_data = 16'b1000011010111100;
    else if (pixel_index == 4483) oled_data = 16'b0110111001111010;
    else if (pixel_index == 4495) oled_data = 16'b0110111010111101;
    else if (pixel_index == 4502 || pixel_index == 4505) oled_data = 16'b0101111011111101;
    else if (pixel_index == 4511) oled_data = 16'b0110111011111100;
    else if (pixel_index == 4512 || pixel_index == 5425) oled_data = 16'b0010100110001000;
    else if (pixel_index == 4514) oled_data = 16'b0010000110001001;
    else if (pixel_index == 4515) oled_data = 16'b0010100101001000;
    else if (pixel_index == 4516) oled_data = 16'b0010000111001010;
    else if (pixel_index == 4517) oled_data = 16'b0010101001001011;
    else if (pixel_index == 4518) oled_data = 16'b0011001000001101;
    else if (pixel_index == 4519) oled_data = 16'b0011001000001100;
    else if (pixel_index == 4520) oled_data = 16'b0011101001001011;
    else if (pixel_index == 4521 || pixel_index == 6063) oled_data = 16'b0011101010001100;
    else if (pixel_index == 4522 || pixel_index == 5250 || pixel_index == 5367) oled_data = 16'b0100001010001100;
    else if (pixel_index == 4523 || pixel_index == 5372 || pixel_index == 6082) oled_data = 16'b0011001000001011;
    else if (pixel_index == 4524) oled_data = 16'b0100001000001100;
    else if (pixel_index == 4525 || pixel_index == 6006) oled_data = 16'b0011101000001100;
    else if (pixel_index == 4526 || ((pixel_index >= 5373) && (pixel_index <= 5374)) || pixel_index == 5980) oled_data = 16'b0100001001001100;
    else if (pixel_index == 4527 || pixel_index == 5162 || pixel_index == 5173) oled_data = 16'b0100001011001111;
    else if (pixel_index == 4528) oled_data = 16'b0101001100010000;
    else if (pixel_index == 4529) oled_data = 16'b0101101101010000;
    else if (pixel_index == 4532 || pixel_index == 4620 || pixel_index == 4623 || ((pixel_index >= 5181) && (pixel_index <= 5182)) || pixel_index == 5895 || pixel_index == 5967) oled_data = 16'b0111110000010010;
    else if (pixel_index == 4533 || pixel_index == 4617 || pixel_index == 4624 || pixel_index == 4706 || pixel_index == 5274) oled_data = 16'b0111110001010011;
    else if (pixel_index == 4534 || pixel_index == 4900 || pixel_index == 5001 || (pixel_index >= 5275) && (pixel_index <= 5276)) oled_data = 16'b1000010001010011;
    else if (pixel_index == 4535) oled_data = 16'b1000010011110101;
    else if (pixel_index == 4536 || pixel_index == 4986) oled_data = 16'b1001010011110110;
    else if (pixel_index == 4537 || pixel_index == 4800 || pixel_index == 4902 || pixel_index == 4983 || pixel_index == 5128 || pixel_index == 5433 || pixel_index == 6126) oled_data = 16'b1010110110110111;
    else if (pixel_index == 4539 || pixel_index == 4978 || pixel_index == 5006 || pixel_index == 5235) oled_data = 16'b1011010111111000;
    else if (pixel_index == 4540 || pixel_index == 4985 || pixel_index == 5617 || pixel_index == 5760) oled_data = 16'b1100011000111001;
    else if (pixel_index == 4542 || pixel_index == 4632 || pixel_index == 5126 || pixel_index == 5465) oled_data = 16'b1100011000111010;
    else if (((pixel_index >= 4543) && (pixel_index <= 4544)) || pixel_index == 4684 || pixel_index == 4686 || pixel_index == 4912 || pixel_index == 5234 || pixel_index == 5356) oled_data = 16'b1100111010111011;
    else if (pixel_index == 4551 || pixel_index == 4699 || pixel_index == 4701 || pixel_index == 4878) oled_data = 16'b1100011010111100;
    else if (pixel_index == 4552) oled_data = 16'b1100011011111011;
    else if (pixel_index == 4554) oled_data = 16'b1010011001111001;
    else if (pixel_index == 4556) oled_data = 16'b1011011001111011;
    else if (pixel_index == 4557 || pixel_index == 5790) oled_data = 16'b1000110000010001;
    else if (pixel_index == 4558) oled_data = 16'b0101101000001010;
    else if (pixel_index == 4560 || pixel_index == 5956) oled_data = 16'b0110001110001111;
    else if (pixel_index == 4589) oled_data = 16'b1001011001111010;
    else if (pixel_index == 4591) oled_data = 16'b1010111011111100;
    else if (pixel_index == 4598) oled_data = 16'b1001111011111100;
    else if (pixel_index == 4608) oled_data = 16'b0100101100001110;
    else if (pixel_index == 4610 || pixel_index == 5158 || pixel_index == 5257) oled_data = 16'b0101001100001111;
    else if (pixel_index == 4611) oled_data = 16'b0101101011001110;
    else if (pixel_index == 4612 || pixel_index == 5177) oled_data = 16'b0101101100010000;
    else if (pixel_index == 4615 || pixel_index == 5968) oled_data = 16'b0111110000010011;
    else if (pixel_index == 4616) oled_data = 16'b1000010001010100;
    else if (pixel_index == 4618 || pixel_index == 5073 || pixel_index == 5246) oled_data = 16'b1000010000010011;
    else if (pixel_index == 4619) oled_data = 16'b0111010000010011;
    else if (pixel_index == 4622) oled_data = 16'b0111110000010001;
    else if (pixel_index == 4625) oled_data = 16'b0111110001010100;
    else if (pixel_index == 4626 || pixel_index == 5467 || pixel_index == 5806) oled_data = 16'b1001010011110100;
    else if (((pixel_index >= 4627) && (pixel_index <= 4628)) || pixel_index == 4749 || pixel_index == 5468 || pixel_index == 5799) oled_data = 16'b1010010100110101;
    else if (pixel_index == 4629 || pixel_index == 5881 || pixel_index == 5898) oled_data = 16'b1010010101110110;
    else if (pixel_index == 4630 || pixel_index == 4710 || pixel_index == 5807) oled_data = 16'b1010110110110110;
    else if (pixel_index == 4631) oled_data = 16'b1011110111111001;
    else if (pixel_index == 4633 || pixel_index == 4635 || pixel_index == 5695 || pixel_index == 5871 || pixel_index == 6130) oled_data = 16'b1101111010111010;
    else if (pixel_index == 4634 || pixel_index == 5054 || pixel_index == 5377 || pixel_index == 5383 || pixel_index == 5481 || pixel_index == 5525 || pixel_index == 5577 || pixel_index == 5671 || pixel_index == 5673 || pixel_index == 5680 || pixel_index == 5698 || pixel_index == 5702 || pixel_index == 5707 || pixel_index == 6132) oled_data = 16'b1110011011111011;
    else if (pixel_index == 4636 || pixel_index == 4650 || pixel_index == 5124 || pixel_index == 5474 || ((pixel_index >= 5569) && (pixel_index <= 5570)) || pixel_index == 5574 || pixel_index == 5672 || pixel_index == 5693 || pixel_index == 5720 || pixel_index == 5762 || pixel_index == 5768 || ((pixel_index >= 5874) && (pixel_index <= 5875)) || pixel_index == 5921) oled_data = 16'b1101111011111011;
    else if (pixel_index == 4637 || pixel_index == 5227 || pixel_index == 5285 || pixel_index == 5670 || pixel_index == 5675 || pixel_index == 5679 || pixel_index == 5703 || pixel_index == 6114 || (pixel_index >= 6116) && (pixel_index <= 6117)) oled_data = 16'b1110011100111011;
    else if (pixel_index == 4638 || pixel_index == 4667 || pixel_index == 4671 || pixel_index == 4713 || pixel_index == 4891 || pixel_index == 5289 || ((pixel_index >= 5378) && (pixel_index <= 5379)) || ((pixel_index >= 5386) && (pixel_index <= 5387)) || pixel_index == 5566 || ((pixel_index >= 5618) && (pixel_index <= 5619)) || ((pixel_index >= 5676) && (pixel_index <= 5677)) || pixel_index == 5701 || pixel_index == 6000) oled_data = 16'b1101111100111100;
    else if (pixel_index == 4639 || pixel_index == 4652 || pixel_index == 4674 || pixel_index == 4736 || pixel_index == 4876 || pixel_index == 4890 || pixel_index == 4893 || pixel_index == 5012 || pixel_index == 5186 || pixel_index == 5189 || pixel_index == 5286 || pixel_index == 5381 || ((pixel_index >= 5564) && (pixel_index <= 5565)) || pixel_index == 5585 || pixel_index == 5590 || pixel_index == 5660 || pixel_index == 5674 || pixel_index == 5686 || pixel_index == 5691 || ((pixel_index >= 5779) && (pixel_index <= 5781)) || pixel_index == 6031) oled_data = 16'b1110011100111100;
    else if (pixel_index == 4640 || pixel_index == 4977 || pixel_index == 5563 || pixel_index == 5573 || pixel_index == 5669 || pixel_index == 5699 || pixel_index == 5771) oled_data = 16'b1101111100111011;
    else if (pixel_index == 4641 || pixel_index == 4746 || pixel_index == 5296 || ((pixel_index >= 5312) && (pixel_index <= 5313)) || pixel_index == 5552 || pixel_index == 5821) oled_data = 16'b1110011110111101;
    else if (pixel_index == 4642 || ((pixel_index >= 4647) && (pixel_index <= 4648)) || ((pixel_index >= 4733) && (pixel_index <= 4734)) || pixel_index == 4737 || pixel_index == 4744 || pixel_index == 4747 || ((pixel_index >= 4776) && (pixel_index <= 4778)) || pixel_index == 4780 || pixel_index == 4789 || pixel_index == 4874 || pixel_index == 4917 || ((pixel_index >= 4950) && (pixel_index <= 4951)) || pixel_index == 5029 || pixel_index == 5045 || pixel_index == 5305 || pixel_index == 5309 || pixel_index == 5388 || pixel_index == 5390 || pixel_index == 5396 || pixel_index == 5405 || pixel_index == 5460 || pixel_index == 5485 || pixel_index == 5502 || pixel_index == 5562 || pixel_index == 5654 || pixel_index == 5658 || pixel_index == 5716 || pixel_index == 5718 || pixel_index == 5724 || pixel_index == 5852 || pixel_index == 5923 || pixel_index == 6021) oled_data = 16'b1110111101111101;
    else if (pixel_index == 4643 || pixel_index == 4775 || pixel_index == 4822 || pixel_index == 4851 || pixel_index == 4869 || pixel_index == 4948 || pixel_index == 5446 || ((pixel_index >= 5555) && (pixel_index <= 5556)) || pixel_index == 5645 || pixel_index == 5741 || pixel_index == 5826 || (pixel_index >= 6134) && (pixel_index <= 6137)) oled_data = 16'b1111111110111101;
    else if (pixel_index == 4644 || pixel_index == 4755 || pixel_index == 4760 || pixel_index == 4766 || pixel_index == 4770 || pixel_index == 4821 || pixel_index == 4823 || pixel_index == 4838 || pixel_index == 4856 || pixel_index == 4860 || pixel_index == 4867 || pixel_index == 4873 || pixel_index == 4926 || pixel_index == 4937 || pixel_index == 4955 || pixel_index == 5016 || pixel_index == 5021 || pixel_index == 5025 || pixel_index == 5116 || pixel_index == 5204 || pixel_index == 5225 || pixel_index == 5398 || pixel_index == 5445 || pixel_index == 5455 || pixel_index == 5609 || pixel_index == 5632 || pixel_index == 5740 || pixel_index == 5827 || pixel_index == 5834 || pixel_index == 5838 || pixel_index == 5935 || pixel_index == 5943 || pixel_index == 5949 || pixel_index == 6028 || pixel_index == 6042 || pixel_index == 6045) oled_data = 16'b1111111110111110;
    else if (((pixel_index >= 4645) && (pixel_index <= 4646)) || pixel_index == 4651 || pixel_index == 4732 || ((pixel_index >= 4794) && (pixel_index <= 4795)) || ((pixel_index >= 4797) && (pixel_index <= 4798)) || pixel_index == 4854 || pixel_index == 4871 || pixel_index == 4875 || pixel_index == 4887 || ((pixel_index >= 4924) && (pixel_index <= 4925)) || pixel_index == 4947 || pixel_index == 5015 || pixel_index == 5047 || pixel_index == 5050 || pixel_index == 5052 || pixel_index == 5099 || pixel_index == 5122 || pixel_index == 5487 || pixel_index == 5496 || pixel_index == 5531 || pixel_index == 5535 || pixel_index == 5561 || pixel_index == 5601 || pixel_index == 5612 || pixel_index == 5644 || pixel_index == 5650 || pixel_index == 5655 || pixel_index == 6041) oled_data = 16'b1111011101111101;
    else if (pixel_index == 4649 || pixel_index == 4916 || pixel_index == 4953 || pixel_index == 5013 || pixel_index == 5098 || pixel_index == 5190 || pixel_index == 5192 || pixel_index == 5331 || pixel_index == 5484 || pixel_index == 5488 || pixel_index == 5579 || pixel_index == 5595 || pixel_index == 5661 || pixel_index == 5683 || pixel_index == 5685 || pixel_index == 5813 || (pixel_index >= 5822) && (pixel_index <= 5823)) oled_data = 16'b1110111101111100;
    else if (pixel_index == 4653) oled_data = 16'b1010010010110100;
    else if (pixel_index == 4654 || pixel_index == 5134) oled_data = 16'b0111001100001110;
    else if (pixel_index == 4655) oled_data = 16'b0101001001001010;
    else if (pixel_index == 4656) oled_data = 16'b1000110001010000;
    else if (pixel_index == 4657 || pixel_index == 4739 || pixel_index == 4759 || pixel_index == 4791 || pixel_index == 4799 || pixel_index == 4836 || pixel_index == 4866 || pixel_index == 4868 || pixel_index == 4870 || pixel_index == 4872 || pixel_index == 4918 || pixel_index == 4931 || pixel_index == 4952 || pixel_index == 5017 || pixel_index == 5108 || pixel_index == 5191 || pixel_index == 5208 || pixel_index == 5211 || pixel_index == 5301 || pixel_index == 5399 || pixel_index == 5401 || pixel_index == 5452 || pixel_index == 5536 || pixel_index == 5554 || pixel_index == 5607 || pixel_index == 5620 || pixel_index == 5624 || pixel_index == 5647 || ((pixel_index >= 5651) && (pixel_index <= 5652)) || pixel_index == 5743 || ((pixel_index >= 5747) && (pixel_index <= 5750)) || pixel_index == 5756 || pixel_index == 5825 || pixel_index == 5853 || pixel_index == 5926 || pixel_index == 5929 || pixel_index == 5931 || pixel_index == 6025 || pixel_index == 6029) oled_data = 16'b1111011110111101;
    else if (pixel_index == 4658 || pixel_index == 4735 || pixel_index == 4765 || pixel_index == 4930 || pixel_index == 5028 || ((pixel_index >= 5030) && (pixel_index <= 5031)) || pixel_index == 5111 || pixel_index == 5195 || pixel_index == 5287 || pixel_index == 5300 || pixel_index == 5303 || pixel_index == 5406 || pixel_index == 5494 || pixel_index == 5504 || pixel_index == 5509 || pixel_index == 5547 || pixel_index == 5605 || pixel_index == 5610 || ((pixel_index >= 5656) && (pixel_index <= 5657)) || pixel_index == 5689 || pixel_index == 5925 || pixel_index == 6023) oled_data = 16'b1110111101111110;
    else if (pixel_index == 4659 || pixel_index == 4885 || pixel_index == 5033 || ((pixel_index >= 5095) && (pixel_index <= 5096)) || pixel_index == 5376 || pixel_index == 5395 || pixel_index == 5417 || pixel_index == 5479 || pixel_index == 5592 || pixel_index == 5684 || pixel_index == 5687 || pixel_index == 5819) oled_data = 16'b1110011100111101;
    else if (pixel_index == 4660) oled_data = 16'b1101111101111110;
    else if (pixel_index == 4663 || pixel_index == 5043 || pixel_index == 5206 || pixel_index == 5281) oled_data = 16'b1101111101111101;
    else if (pixel_index == 4665 || pixel_index == 5473 || pixel_index == 5665) oled_data = 16'b1101111010111100;
    else if (pixel_index == 4668 || pixel_index == 4675 || pixel_index == 4895 || pixel_index == 5094 || pixel_index == 5480 || pixel_index == 5568 || ((pixel_index >= 5575) && (pixel_index <= 5576)) || pixel_index == 5666 || pixel_index == 5694 || pixel_index == 5767 || pixel_index == 5770 || pixel_index == 6118) oled_data = 16'b1101111011111100;
    else if (pixel_index == 4670 || pixel_index == 4680 || pixel_index == 4884 || pixel_index == 4913 || pixel_index == 5571 || (pixel_index >= 6119) && (pixel_index <= 6120)) oled_data = 16'b1101111011111101;
    else if (pixel_index == 4672) oled_data = 16'b1101011100111101;
    else if (pixel_index == 4677 || pixel_index == 4691 || pixel_index == 4975) oled_data = 16'b1100111011111011;
    else if (pixel_index == 4683 || pixel_index == 5332 || pixel_index == 5354 || pixel_index == 5667 || pixel_index == 5714 || pixel_index == 5999 || pixel_index == 6129) oled_data = 16'b1101011011111100;
    else if (pixel_index == 4690) oled_data = 16'b1100111100111100;
    else if (pixel_index == 4704) oled_data = 16'b0111010001010010;
    else if (pixel_index == 4708) oled_data = 16'b1000110001010100;
    else if (pixel_index == 4709 || pixel_index == 5057 || pixel_index == 5062) oled_data = 16'b1001110011110101;
    else if (pixel_index == 4711 || pixel_index == 5522 || pixel_index == 5814) oled_data = 16'b1011111000110111;
    else if (pixel_index == 4712 || pixel_index == 5140) oled_data = 16'b1100011001111000;
    else if (((pixel_index >= 4714) && (pixel_index <= 4715)) || pixel_index == 4743 || pixel_index == 4787 || pixel_index == 4796 || pixel_index == 4808 || pixel_index == 4886 || pixel_index == 4915 || pixel_index == 5044 || pixel_index == 5290 || pixel_index == 5393 || pixel_index == 5482 || pixel_index == 5583 || ((pixel_index >= 5586) && (pixel_index <= 5588)) || pixel_index == 5600 || pixel_index == 5662 || pixel_index == 5690 || pixel_index == 5811 || pixel_index == 6022) oled_data = 16'b1110111100111101;
    else if (pixel_index == 4716 || pixel_index == 5199 || pixel_index == 5397 || pixel_index == 5409 || pixel_index == 5415 || pixel_index == 5511 || pixel_index == 5545 || pixel_index == 5649 || pixel_index == 5730 || pixel_index == 5828 || pixel_index == 5940) oled_data = 16'b1111011101111111;
    else if (pixel_index == 4717 || pixel_index == 4783 || pixel_index == 4809 || pixel_index == 4815 || ((pixel_index >= 4852) && (pixel_index <= 4853)) || pixel_index == 4921 || pixel_index == 5023 || pixel_index == 5027 || pixel_index == 5207 || pixel_index == 5222 || pixel_index == 5295 || pixel_index == 5297 || ((pixel_index >= 5306) && (pixel_index <= 5307)) || pixel_index == 5413 || pixel_index == 5495 || pixel_index == 5507 || pixel_index == 5604 || pixel_index == 5606 || pixel_index == 5726 || ((pixel_index >= 5744) && (pixel_index <= 5746)) || pixel_index == 5759 || pixel_index == 5812 || pixel_index == 5841 || pixel_index == 5905 || pixel_index == 5934 || pixel_index == 6026) oled_data = 16'b1110111110111110;
    else if (((pixel_index >= 4718) && (pixel_index <= 4719)) || ((pixel_index >= 4763) && (pixel_index <= 4764)) || pixel_index == 4773 || pixel_index == 4793 || pixel_index == 4830 || pixel_index == 4850 || pixel_index == 4923 || pixel_index == 5051 || ((pixel_index >= 5292) && (pixel_index <= 5293)) || pixel_index == 5314 || pixel_index == 5486 || pixel_index == 5497 || pixel_index == 5548 || pixel_index == 5629 || pixel_index == 5638 || pixel_index == 5734 || pixel_index == 5758 || pixel_index == 5833 || pixel_index == 5904 || pixel_index == 5924 || pixel_index == 6027) oled_data = 16'b1111011101111110;
    else if (pixel_index == 4720 || pixel_index == 4738 || pixel_index == 4756 || pixel_index == 4768 || pixel_index == 4771 || pixel_index == 4786 || pixel_index == 4790 || pixel_index == 4792 || ((pixel_index >= 4810) && (pixel_index <= 4811)) || pixel_index == 4814 || pixel_index == 4817 || pixel_index == 4819 || ((pixel_index >= 4827) && (pixel_index <= 4829)) || ((pixel_index >= 4831) && (pixel_index <= 4832)) || pixel_index == 4837 || pixel_index == 4839 || pixel_index == 4855 || ((pixel_index >= 4881) && (pixel_index <= 4882)) || pixel_index == 4888 || pixel_index == 4932 || pixel_index == 5196 || pixel_index == 5209 || pixel_index == 5216 || pixel_index == 5218 || pixel_index == 5223 || ((pixel_index >= 5298) && (pixel_index <= 5299)) || pixel_index == 5304 || pixel_index == 5319 || pixel_index == 5404 || pixel_index == 5414 || pixel_index == 5456 || pixel_index == 5501 || ((pixel_index >= 5539) && (pixel_index <= 5540)) || pixel_index == 5608 || pixel_index == 5627 || pixel_index == 5631 || pixel_index == 5634 || pixel_index == 5637 || pixel_index == 5643 || pixel_index == 5721 || pixel_index == 5723 || pixel_index == 5729 || pixel_index == 5733 || pixel_index == 5738 || pixel_index == 5751 || ((pixel_index >= 5753) && (pixel_index <= 5755)) || pixel_index == 5757 || ((pixel_index >= 5830) && (pixel_index <= 5832)) || pixel_index == 5835 || pixel_index == 5851 || pixel_index == 5854 || pixel_index == 5933 || pixel_index == 5944 || ((pixel_index >= 5947) && (pixel_index <= 5948)) || pixel_index == 6040 || pixel_index == 6138) oled_data = 16'b1111011110111110;
    else if (pixel_index == 4721 || pixel_index == 4723 || pixel_index == 4731 || pixel_index == 4785 || pixel_index == 4813 || pixel_index == 4861 || pixel_index == 4880 || pixel_index == 4920 || pixel_index == 5107 || ((pixel_index >= 5117) && (pixel_index <= 5118)) || pixel_index == 5202 || pixel_index == 5213 || pixel_index == 5450 || pixel_index == 5551 || pixel_index == 5839 || pixel_index == 5843 || ((pixel_index >= 5846) && (pixel_index <= 5847)) || pixel_index == 5927 || pixel_index == 5937 || pixel_index == 5942 || pixel_index == 6046) oled_data = 16'b1111011111111110;
    else if (pixel_index == 4722 || pixel_index == 4927 || pixel_index == 4936 || pixel_index == 5018 || pixel_index == 5022 || pixel_index == 5101 || pixel_index == 5459 || pixel_index == 5541 || pixel_index == 5544 || pixel_index == 5621 || pixel_index == 5625 || pixel_index == 5829 || pixel_index == 5844 || pixel_index == 5928 || pixel_index == 5939 || pixel_index == 6039) oled_data = 16'b1111111110111111;
    else if (((pixel_index >= 4724) && (pixel_index <= 4725)) || ((pixel_index >= 4729) && (pixel_index <= 4730)) || pixel_index == 4761 || pixel_index == 4812 || pixel_index == 4933 || pixel_index == 4935 || pixel_index == 5020 || pixel_index == 5024 || ((pixel_index >= 5105) && (pixel_index <= 5106)) || pixel_index == 5203 || pixel_index == 5311 || pixel_index == 5317 || ((pixel_index >= 5320) && (pixel_index <= 5321)) || pixel_index == 5447 || pixel_index == 5449 || ((pixel_index >= 5457) && (pixel_index <= 5458)) || pixel_index == 5532 || pixel_index == 5538 || pixel_index == 5543 || pixel_index == 5622 || pixel_index == 5626 || pixel_index == 5636 || pixel_index == 5945 || pixel_index == 6043) oled_data = 16'b1111111111111111;
    else if (pixel_index == 4726 || pixel_index == 4842 || pixel_index == 4849 || pixel_index == 5103 || pixel_index == 5224 || ((pixel_index >= 5410) && (pixel_index <= 5412)) || pixel_index == 5500 || pixel_index == 5623) oled_data = 16'b1111011111111101;
    else if (((pixel_index >= 4727) && (pixel_index <= 4728)) || pixel_index == 4754 || pixel_index == 4820 || pixel_index == 4835 || pixel_index == 4841 || pixel_index == 4859 || pixel_index == 4862 || pixel_index == 4865 || pixel_index == 4928 || ((pixel_index >= 4938) && (pixel_index <= 4939)) || pixel_index == 5019 || pixel_index == 5210 || pixel_index == 5212 || pixel_index == 5217 || pixel_index == 5316 || pixel_index == 5318 || pixel_index == 5451 || pixel_index == 5498 || pixel_index == 5534 || pixel_index == 5542 || pixel_index == 5633 || pixel_index == 5717 || ((pixel_index >= 5727) && (pixel_index <= 5728)) || pixel_index == 5737 || pixel_index == 5845 || pixel_index == 5936 || ((pixel_index >= 5950) && (pixel_index <= 5951)) || pixel_index == 6044 || pixel_index == 6047) oled_data = 16'b1111111111111110;
    else if (pixel_index == 4740 || pixel_index == 5110 || pixel_index == 5121 || pixel_index == 5194 || pixel_index == 5198 || pixel_index == 5330 || pixel_index == 5490 || pixel_index == 5611 || pixel_index == 5646 || pixel_index == 6133) oled_data = 16'b1111011101111100;
    else if (pixel_index == 4741 || pixel_index == 4889 || pixel_index == 5408 || pixel_index == 5499 || pixel_index == 5512 || pixel_index == 5855 || pixel_index == 6032 || pixel_index == 6034) oled_data = 16'b1111111101111101;
    else if (pixel_index == 4742 || pixel_index == 4772 || pixel_index == 5014 || pixel_index == 5193 || pixel_index == 5560) oled_data = 16'b1111011100111101;
    else if (pixel_index == 4748 || pixel_index == 5580) oled_data = 16'b1110011101111011;
    else if (pixel_index == 4751) oled_data = 16'b0101101001001010;
    else if (pixel_index == 4752 || pixel_index == 5325) oled_data = 16'b0111101101001111;
    else if (pixel_index == 4753 || ((pixel_index >= 4824) && (pixel_index <= 4825)) || pixel_index == 4863 || pixel_index == 4934 || pixel_index == 5100 || pixel_index == 5104 || pixel_index == 5448 || pixel_index == 5630 || pixel_index == 5635 || ((pixel_index >= 5639) && (pixel_index <= 5640)) || ((pixel_index >= 5735) && (pixel_index <= 5736)) || pixel_index == 5842 || pixel_index == 5850 || pixel_index == 5946 || pixel_index == 6037) oled_data = 16'b1111011111111111;
    else if (pixel_index == 4757 || pixel_index == 4788 || pixel_index == 5493 || pixel_index == 5553 || pixel_index == 5589 || pixel_index == 5594 || pixel_index == 5596 || pixel_index == 5678 || pixel_index == 5688 || pixel_index == 5922 || pixel_index == 6030) oled_data = 16'b1110011101111101;
    else if (pixel_index == 4758 || pixel_index == 5291 || pixel_index == 5392 || pixel_index == 5489 || pixel_index == 5505 || pixel_index == 5559 || pixel_index == 5578 || pixel_index == 5584 || pixel_index == 5598 || pixel_index == 5613 || pixel_index == 5615 || pixel_index == 5659 || pixel_index == 5682 || pixel_index == 5818 || pixel_index == 5824) oled_data = 16'b1110111100111100;
    else if (pixel_index == 4762 || pixel_index == 5109 || pixel_index == 5530 || pixel_index == 5550 || pixel_index == 5602 || pixel_index == 5906) oled_data = 16'b1111011110111100;
    else if (pixel_index == 4767 || pixel_index == 5528 || pixel_index == 6142) oled_data = 16'b1110011110111111;
    else if (pixel_index == 4769 || pixel_index == 4919 || pixel_index == 5840 || pixel_index == 5848) oled_data = 16'b1110111111111110;
    else if (pixel_index == 4774 || pixel_index == 5200 || pixel_index == 5315) oled_data = 16'b1111111101111110;
    else if (pixel_index == 4779 || pixel_index == 4781 || pixel_index == 5454 || pixel_index == 5603 || pixel_index == 5628 || pixel_index == 5653 || pixel_index == 6019) oled_data = 16'b1110111110111100;
    else if (pixel_index == 4784 || pixel_index == 4826 || ((pixel_index >= 4833) && (pixel_index <= 4834)) || pixel_index == 4840 || pixel_index == 4858 || pixel_index == 4864 || pixel_index == 4929 || pixel_index == 4954 || pixel_index == 5026 || pixel_index == 5205 || pixel_index == 5219 || pixel_index == 5310 || pixel_index == 5403 || ((pixel_index >= 5442) && (pixel_index <= 5444)) || pixel_index == 5508 || pixel_index == 5510 || pixel_index == 5529 || pixel_index == 5641 || pixel_index == 5648 || pixel_index == 5722 || ((pixel_index >= 5731) && (pixel_index <= 5732)) || pixel_index == 5739 || pixel_index == 5752 || ((pixel_index >= 5836) && (pixel_index <= 5837)) || pixel_index == 5849 || pixel_index == 5932 || pixel_index == 5938 || pixel_index == 5941 || pixel_index == 6024 || pixel_index == 6038 || pixel_index == 6139) oled_data = 16'b1111011110111111;
    else if (pixel_index == 4801 || pixel_index == 5323 || pixel_index == 6127) oled_data = 16'b1011010110110111;
    else if (pixel_index == 4802) oled_data = 16'b1011011000111000;
    else if (((pixel_index >= 4803) && (pixel_index <= 4804)) || pixel_index == 5131 || pixel_index == 5865) oled_data = 16'b1100011000111000;
    else if (pixel_index == 4805 || pixel_index == 4908 || pixel_index == 4911 || pixel_index == 4960 || pixel_index == 5008 || pixel_index == 5185 || pixel_index == 5333 || ((pixel_index >= 5352) && (pixel_index <= 5353)) || pixel_index == 5664 || pixel_index == 5915) oled_data = 16'b1100111001111010;
    else if (pixel_index == 4806 || pixel_index == 5706 || pixel_index == 5708 || pixel_index == 5769 || pixel_index == 5876 || pixel_index == 5903) oled_data = 16'b1101111010111011;
    else if (pixel_index == 4816 || pixel_index == 4922 || pixel_index == 5046 || pixel_index == 5102 || pixel_index == 5226 || pixel_index == 5537 || pixel_index == 5642 || (pixel_index >= 6140) && (pixel_index <= 6141)) oled_data = 16'b1110111110111111;
    else if (pixel_index == 4818 || pixel_index == 5115 || pixel_index == 5201) oled_data = 16'b1111111101111111;
    else if (pixel_index == 4844 || pixel_index == 4892 || pixel_index == 5355 || pixel_index == 5476 || pixel_index == 5567 || pixel_index == 5668 || pixel_index == 5772) oled_data = 16'b1101011011111011;
    else if (pixel_index == 4845 || pixel_index == 5247) oled_data = 16'b1001110010110100;
    else if (pixel_index == 4846 || pixel_index == 6048) oled_data = 16'b0111101110001111;
    else if (pixel_index == 4847) oled_data = 16'b0110001010001100;
    else if (pixel_index == 4848) oled_data = 16'b1000001111001111;
    else if (pixel_index == 4857 || pixel_index == 4949 || pixel_index == 5214 || pixel_index == 5402 || pixel_index == 5930) oled_data = 16'b1111111111111101;
    else if (pixel_index == 4879 || pixel_index == 5032 || pixel_index == 5503 || pixel_index == 5527) oled_data = 16'b1110011101111110;
    else if (pixel_index == 4883) oled_data = 16'b1110011011111101;
    else if (pixel_index == 4896 || pixel_index == 5979) oled_data = 16'b0101001011001110;
    else if (pixel_index == 4897 || pixel_index == 5885) oled_data = 16'b0101101011001101;
    else if (pixel_index == 4898 || pixel_index == 6100) oled_data = 16'b0111001110001111;
    else if (pixel_index == 4901 || pixel_index == 5060) oled_data = 16'b1001010010110101;
    else if (pixel_index == 4903 || pixel_index == 5055) oled_data = 16'b1011111001111001;
    else if (pixel_index == 4904 || pixel_index == 4962 || pixel_index == 5093 || pixel_index == 5125 || pixel_index == 6128) oled_data = 16'b1100011001111010;
    else if (pixel_index == 4905 || pixel_index == 5138) oled_data = 16'b1100010111111010;
    else if (pixel_index == 4906 || pixel_index == 5141) oled_data = 16'b1011111000111010;
    else if (pixel_index == 4907 || pixel_index == 4961) oled_data = 16'b1100111000111010;
    else if (pixel_index == 4909 || pixel_index == 5783) oled_data = 16'b1101111011111001;
    else if (pixel_index == 4910) oled_data = 16'b1100111011111001;
    else if (pixel_index == 4914 || pixel_index == 5817) oled_data = 16'b1110011010111100;
    else if (pixel_index == 4940) oled_data = 16'b1100011000111011;
    else if (pixel_index == 4941 || pixel_index == 5789) oled_data = 16'b1000110000010011;
    else if (pixel_index == 4942 || pixel_index == 5963) oled_data = 16'b0111001111001111;
    else if (pixel_index == 4943 || pixel_index == 5230 || pixel_index == 6055 || pixel_index == 6062) oled_data = 16'b0101001010001100;
    else if (pixel_index == 4944) oled_data = 16'b1000101110001110;
    else if (pixel_index == 4945) oled_data = 16'b1111111111111011;
    else if (pixel_index == 4946 || pixel_index == 4956 || (pixel_index >= 5119) && (pixel_index <= 5120)) oled_data = 16'b1110011110111110;
    else if (pixel_index == 4958 || pixel_index == 5436 || pixel_index == 5873) oled_data = 16'b1101011010111011;
    else if (pixel_index == 4959) oled_data = 16'b1100110111111001;
    else if (((pixel_index >= 4964) && (pixel_index <= 4965)) || pixel_index == 5742) oled_data = 16'b1111111110111100;
    else if (pixel_index == 4966) oled_data = 16'b1111111110111011;
    else if (pixel_index == 4967 || pixel_index == 4969 || pixel_index == 4976) oled_data = 16'b1111011110111011;
    else if (pixel_index == 4968) oled_data = 16'b1111111111111100;
    else if (pixel_index == 4970) oled_data = 16'b1110111101111010;
    else if (pixel_index == 4971 || pixel_index == 5437) oled_data = 16'b1101011011111010;
    else if (pixel_index == 4972 || pixel_index == 5359) oled_data = 16'b1010110110111001;
    else if (pixel_index == 4973) oled_data = 16'b0111010010111001;
    else if (pixel_index == 4974) oled_data = 16'b0110010000011010;
    else if (pixel_index == 4979) oled_data = 16'b1000010001010110;
    else if (pixel_index == 4980) oled_data = 16'b0110001110010101;
    else if (pixel_index == 4981) oled_data = 16'b0111110000010101;
    else if (pixel_index == 4982 || pixel_index == 5005) oled_data = 16'b1010110101110111;
    else if (pixel_index == 4984 || pixel_index == 5036 || pixel_index == 5127 || pixel_index == 5358 || pixel_index == 5808 || pixel_index == 5861) oled_data = 16'b1011110111111000;
    else if (pixel_index == 4987 || pixel_index == 4990) oled_data = 16'b1000010010110101;
    else if (pixel_index == 4989) oled_data = 16'b0111110010110101;
    else if (pixel_index == 4991) oled_data = 16'b0111010001010101;
    else if (pixel_index == 4992) oled_data = 16'b0100101001001011;
    else if (pixel_index == 4993 || pixel_index == 5231 || pixel_index == 5252) oled_data = 16'b0100001001001011;
    else if (pixel_index == 4994 || pixel_index == 6053) oled_data = 16'b0101101100001110;
    else if (pixel_index == 4998 || pixel_index == 5977) oled_data = 16'b0110101101001111;
    else if (pixel_index == 4999 || pixel_index == 5153) oled_data = 16'b0111001110010000;
    else if (pixel_index == 5000 || pixel_index == 5975) oled_data = 16'b0111101111010001;
    else if (pixel_index == 5002 || pixel_index == 5065) oled_data = 16'b1000010010110100;
    else if (pixel_index == 5003) oled_data = 16'b1000110010110101;
    else if (pixel_index == 5004) oled_data = 16'b1001110101110110;
    else if (pixel_index == 5007 || pixel_index == 5786 || pixel_index == 6089) oled_data = 16'b1011111000111000;
    else if (pixel_index == 5035 || pixel_index == 5384 || pixel_index == 5705 || pixel_index == 5719 || pixel_index == 5763 || pixel_index == 5877 || pixel_index == 6094) oled_data = 16'b1101111011111010;
    else if (pixel_index == 5037) oled_data = 16'b1000101111010000;
    else if (pixel_index == 5038) oled_data = 16'b0110101100001101;
    else if (pixel_index == 5039) oled_data = 16'b0101101001001011;
    else if (pixel_index == 5040) oled_data = 16'b0110101110001110;
    else if (pixel_index == 5041 || pixel_index == 5048 || pixel_index == 5282 || pixel_index == 5513 || pixel_index == 5663 || pixel_index == 5681 || pixel_index == 5692 || pixel_index == 5715 || pixel_index == 6018) oled_data = 16'b1110011011111100;
    else if (pixel_index == 5042 || pixel_index == 5284 || pixel_index == 6131) oled_data = 16'b1110111100111011;
    else if (pixel_index == 5049) oled_data = 16'b1101011110111101;
    else if (pixel_index == 5053 || pixel_index == 5558) oled_data = 16'b1111011100111100;
    else if (pixel_index == 5058) oled_data = 16'b1001010010110100;
    else if (pixel_index == 5059 || pixel_index == 5432) oled_data = 16'b1001110010110101;
    else if (pixel_index == 5061) oled_data = 16'b1001010010110110;
    else if (pixel_index == 5063) oled_data = 16'b1010010100110100;
    else if (pixel_index == 5066 || pixel_index == 5245 || pixel_index == 5279 || pixel_index == 6003 || pixel_index == 6096) oled_data = 16'b1000110011110100;
    else if (pixel_index == 5067) oled_data = 16'b0111110000010100;
    else if (pixel_index == 5068) oled_data = 16'b0110101110010011;
    else if (pixel_index == 5069) oled_data = 16'b0100101011010010;
    else if (pixel_index == 5070) oled_data = 16'b0101001100010010;
    else if (pixel_index == 5071) oled_data = 16'b1001010100110101;
    else if (pixel_index == 5072 || pixel_index == 5470 || pixel_index == 5798) oled_data = 16'b1001110011110100;
    else if (pixel_index == 5074 || pixel_index == 6101) oled_data = 16'b0110101110010010;
    else if (pixel_index == 5075 || pixel_index == 5086) oled_data = 16'b0100101101010001;
    else if (pixel_index == 5076) oled_data = 16'b0100001100010010;
    else if (pixel_index == 5077) oled_data = 16'b0100101101010010;
    else if (pixel_index == 5079) oled_data = 16'b0101101110010010;
    else if (pixel_index == 5081) oled_data = 16'b0110001111010011;
    else if (pixel_index == 5082) oled_data = 16'b0101001101010010;
    else if (pixel_index == 5083 || pixel_index == 5085 || pixel_index == 5087) oled_data = 16'b0100101100010001;
    else if (pixel_index == 5084) oled_data = 16'b0100001011010001;
    else if (pixel_index == 5088 || pixel_index == 5132 || pixel_index == 5787 || pixel_index == 5802) oled_data = 16'b1011010101110110;
    else if (pixel_index == 5090 || pixel_index == 5345 || pixel_index == 5857) oled_data = 16'b1011111000111001;
    else if (pixel_index == 5091) oled_data = 16'b1011110110111010;
    else if (pixel_index == 5092 || pixel_index == 5344 || pixel_index == 5899) oled_data = 16'b1011010110111001;
    else if (pixel_index == 5112 || pixel_index == 5416 || pixel_index == 5441) oled_data = 16'b1110111100111110;
    else if (pixel_index == 5113 || pixel_index == 5407) oled_data = 16'b1111011100111110;
    else if (pixel_index == 5114 || pixel_index == 5215 || pixel_index == 5220 || pixel_index == 5546) oled_data = 16'b1110111101111111;
    else if (pixel_index == 5130 || pixel_index == 5913) oled_data = 16'b1011010111111001;
    else if (pixel_index == 5133) oled_data = 16'b1001010001010001;
    else if (pixel_index == 5136) oled_data = 16'b0100101001001001;
    else if (pixel_index == 5137 || pixel_index == 5816) oled_data = 16'b1011110110111000;
    else if (pixel_index == 5142 || pixel_index == 5709) oled_data = 16'b1101011001111010;
    else if (pixel_index == 5143) oled_data = 16'b1100111000110110;
    else if (pixel_index == 5144 || pixel_index == 5148) oled_data = 16'b1010110011110011;
    else if (pixel_index == 5145 || pixel_index == 5149) oled_data = 16'b1001110010110010;
    else if (pixel_index == 5146) oled_data = 16'b1011010110110101;
    else if (pixel_index == 5147) oled_data = 16'b1100111000110111;
    else if (pixel_index == 5150 || pixel_index == 5953) oled_data = 16'b1001110100110011;
    else if (pixel_index == 5152 || pixel_index == 5971 || pixel_index == 5973) oled_data = 16'b1001010010110010;
    else if (pixel_index == 5154) oled_data = 16'b0110001100001111;
    else if (pixel_index == 5155) oled_data = 16'b0101101011001111;
    else if (pixel_index == 5156 || pixel_index == 5254) oled_data = 16'b0100101010001110;
    else if (pixel_index == 5157 || pixel_index == 5892) oled_data = 16'b0101001010001110;
    else if (pixel_index == 5159 || pixel_index == 5263) oled_data = 16'b0100001010001101;
    else if (pixel_index == 5160) oled_data = 16'b0011101010001110;
    else if (pixel_index == 5161 || ((pixel_index >= 5169) && (pixel_index <= 5170)) || pixel_index == 5174) oled_data = 16'b0011101010001111;
    else if (pixel_index == 5163) oled_data = 16'b0100001011010000;
    else if ((pixel_index >= 5165) && (pixel_index <= 5166)) oled_data = 16'b0101001100001110;
    else if (pixel_index == 5168) oled_data = 16'b0011101001010000;
    else if (pixel_index == 5172) oled_data = 16'b0100101101010000;
    else if (pixel_index == 5175) oled_data = 16'b0100001010010000;
    else if (pixel_index == 5178) oled_data = 16'b0110001101010000;
    else if (((pixel_index >= 5179) && (pixel_index <= 5180)) || pixel_index == 5267) oled_data = 16'b0110101111010001;
    else if (pixel_index == 5183 || pixel_index == 5969) oled_data = 16'b1000010010110011;
    else if (pixel_index == 5184 || pixel_index == 5357) oled_data = 16'b1100010111111001;
    else if (pixel_index == 5221) oled_data = 16'b1101111110111111;
    else if (pixel_index == 5228) oled_data = 16'b1011110101110011;
    else if (pixel_index == 5229) oled_data = 16'b1000010000001110;
    else if (pixel_index == 5232) oled_data = 16'b0010100100000100;
    else if (pixel_index == 5233 || pixel_index == 5788 || pixel_index == 6011) oled_data = 16'b1001110011110011;
    else if (pixel_index == 5236) oled_data = 16'b1010110101111000;
    else if (pixel_index == 5237) oled_data = 16'b1011110101110111;
    else if (pixel_index == 5238) oled_data = 16'b1100010101110111;
    else if (pixel_index == 5239) oled_data = 16'b1001101101001101;
    else if (pixel_index == 5240) oled_data = 16'b0101101010000101;
    else if (pixel_index == 5241) oled_data = 16'b0100000101000001;
    else if (pixel_index == 5242) oled_data = 16'b0101101010001010;
    else if (pixel_index == 5243) oled_data = 16'b1011110110110111;
    else if (pixel_index == 5244 || pixel_index == 5801 || pixel_index == 5901) oled_data = 16'b1010110101110110;
    else if (pixel_index == 5248) oled_data = 16'b1000110000010000;
    else if (pixel_index == 5249) oled_data = 16'b0101101011001010;
    else if (pixel_index == 5253) oled_data = 16'b0101001011001111;
    else if (pixel_index == 5255) oled_data = 16'b0011001000001110;
    else if (pixel_index == 5256) oled_data = 16'b0011101001001110;
    else if (pixel_index == 5258) oled_data = 16'b0100101001001101;
    else if (pixel_index == 5259) oled_data = 16'b0100101001001100;
    else if (pixel_index == 5260) oled_data = 16'b0100001001001101;
    else if (pixel_index == 5261 || pixel_index == 5982 || pixel_index == 5984 || pixel_index == 6068 || pixel_index == 6075 || pixel_index == 6077) oled_data = 16'b0011001000001010;
    else if (pixel_index == 5262) oled_data = 16'b0010100111001011;
    else if ((pixel_index >= 5265) && (pixel_index <= 5266)) oled_data = 16'b0110001110010010;
    else if (pixel_index == 5268) oled_data = 16'b0110001011001110;
    else if ((pixel_index >= 5269) && (pixel_index <= 5270)) oled_data = 16'b0110001011001101;
    else if (pixel_index == 5271 || pixel_index == 6099) oled_data = 16'b0110001101001101;
    else if (pixel_index == 5272 || pixel_index == 6087) oled_data = 16'b1000010000010001;
    else if (pixel_index == 5273 || pixel_index == 6105) oled_data = 16'b1000110001010011;
    else if (pixel_index == 5277) oled_data = 16'b1001110100110101;
    else if (pixel_index == 5280 || pixel_index == 5438) oled_data = 16'b1110011110111010;
    else if (pixel_index == 5283) oled_data = 16'b1111011011111101;
    else if (pixel_index == 5322) oled_data = 16'b1111011111111100;
    else if (pixel_index == 5324) oled_data = 16'b1001010000010010;
    else if (pixel_index == 5328) oled_data = 16'b0000100100000100;
    else if (pixel_index == 5335) oled_data = 16'b1001010011110001;
    else if (pixel_index == 5336) oled_data = 16'b0110101100001011;
    else if (pixel_index == 5337) oled_data = 16'b0100101001001010;
    else if (pixel_index == 5338 || pixel_index == 5990) oled_data = 16'b0101001011001101;
    else if (pixel_index == 5339) oled_data = 16'b1000110010110011;
    else if (pixel_index == 5340) oled_data = 16'b1001110011110110;
    else if (pixel_index == 5341) oled_data = 16'b1001110010110111;
    else if (pixel_index == 5342) oled_data = 16'b1001110011110111;
    else if (pixel_index == 5343) oled_data = 16'b1010010110111000;
    else if (pixel_index == 5346 || pixel_index == 5996 || pixel_index == 6001 || pixel_index == 6110) oled_data = 16'b1100111000111001;
    else if (pixel_index == 5347) oled_data = 16'b1101011001110111;
    else if (pixel_index == 5350) oled_data = 16'b1011011000111011;
    else if (pixel_index == 5360) oled_data = 16'b1100010110111000;
    else if (pixel_index == 5361) oled_data = 16'b1101111000111000;
    else if (pixel_index == 5362 || pixel_index == 5711) oled_data = 16'b1100111001111001;
    else if (pixel_index == 5365) oled_data = 16'b0101101110010000;
    else if (pixel_index == 5366 || pixel_index == 6050) oled_data = 16'b0100101011001110;
    else if (pixel_index == 5368 || pixel_index == 6054) oled_data = 16'b0101001011001100;
    else if (pixel_index == 5369) oled_data = 16'b0101001100001101;
    else if (pixel_index == 5370 || pixel_index == 5375 || pixel_index == 5983 || pixel_index == 6084) oled_data = 16'b0011101000001011;
    else if (pixel_index == 5371) oled_data = 16'b0011000110001010;
    else if (pixel_index == 5382 || pixel_index == 5599 || pixel_index == 5782) oled_data = 16'b1110111011111011;
    else if (pixel_index == 5385 || pixel_index == 5777) oled_data = 16'b1101111100111010;
    else if (pixel_index == 5391 || pixel_index == 5761) oled_data = 16'b1110011011111110;
    else if (pixel_index == 5420) oled_data = 16'b0110001110001100;
    else if (pixel_index == 5421) oled_data = 16'b0101001010001001;
    else if (pixel_index == 5422) oled_data = 16'b0011101000000110;
    else if (pixel_index == 5423) oled_data = 16'b0011100101000101;
    else if (pixel_index == 5424) oled_data = 16'b0010100011000101;
    else if (pixel_index == 5426) oled_data = 16'b0110101110010001;
    else if (pixel_index == 5427 || pixel_index == 5791 || pixel_index == 5952 || pixel_index == 5960) oled_data = 16'b0111101111010000;
    else if (pixel_index == 5428) oled_data = 16'b1001010001010011;
    else if (pixel_index == 5429 || pixel_index == 5471 || pixel_index == 5970) oled_data = 16'b1000110011110011;
    else if (pixel_index == 5430) oled_data = 16'b0111101111010011;
    else if (pixel_index == 5431) oled_data = 16'b1000110010110111;
    else if (pixel_index == 5434) oled_data = 16'b1010111000111001;
    else if (pixel_index == 5435 || pixel_index == 5713) oled_data = 16'b1100111001111011;
    else if (pixel_index == 5439 || pixel_index == 5775) oled_data = 16'b1110111101111011;
    else if (pixel_index == 5440) oled_data = 16'b1110111011111101;
    else if (pixel_index == 5453) oled_data = 16'b1110111111111100;
    else if (pixel_index == 5461 || ((pixel_index >= 5765) && (pixel_index <= 5766)) || pixel_index == 5785 || pixel_index == 5872 || pixel_index == 5917 || pixel_index == 5919 || pixel_index == 6112) oled_data = 16'b1101011010111010;
    else if (pixel_index == 5462) oled_data = 16'b1101111001111010;
    else if (((pixel_index >= 5463) && (pixel_index <= 5464)) || pixel_index == 5809) oled_data = 16'b1101011000111010;
    else if (pixel_index == 5466 || pixel_index == 5469 || pixel_index == 5860) oled_data = 16'b1010110100110110;
    else if (pixel_index == 5472) oled_data = 16'b1110111001111011;
    else if (pixel_index == 5475) oled_data = 16'b1101011100111011;
    else if (pixel_index == 5477) oled_data = 16'b1100111100111011;
    else if (pixel_index == 5483) oled_data = 16'b1110111100111010;
    else if (pixel_index == 5506) oled_data = 16'b1111011101111011;
    else if (pixel_index == 5515) oled_data = 16'b1010110100110011;
    else if (pixel_index == 5517 || pixel_index == 6108) oled_data = 16'b1001010001001111;
    else if (pixel_index == 5519) oled_data = 16'b0101001010001010;
    else if (pixel_index == 5520) oled_data = 16'b0100000111001001;
    else if (pixel_index == 5521) oled_data = 16'b0110101010001111;
    else if (pixel_index == 5526) oled_data = 16'b1111011011111100;
    else if (pixel_index == 5533) oled_data = 16'b1110111111111101;
    else if (pixel_index == 5557) oled_data = 16'b1111011100111011;
    else if (pixel_index == 5572) oled_data = 16'b1101111101111011;
    else if (pixel_index == 5582) oled_data = 16'b1110011101111111;
    else if (pixel_index == 5616) oled_data = 16'b1100111001110111;
    else if (((pixel_index >= 5696) && (pixel_index <= 5697)) || pixel_index == 5920 || pixel_index == 6017 || pixel_index == 6091 || pixel_index == 6115) oled_data = 16'b1110011011111010;
    else if (pixel_index == 5704) oled_data = 16'b1110011010111011;
    else if (pixel_index == 5712) oled_data = 16'b1100111010111000;
    else if (pixel_index == 5764 || pixel_index == 5869 || pixel_index == 6016) oled_data = 16'b1101011001111001;
    else if (pixel_index == 5776 || pixel_index == 5907) oled_data = 16'b1110011100111010;
    else if (pixel_index == 5778) oled_data = 16'b1110111011111100;
    else if (pixel_index == 5784 || pixel_index == 5908 || pixel_index == 5998) oled_data = 16'b1110011010111010;
    else if ((pixel_index >= 5792) && (pixel_index <= 5793)) oled_data = 16'b0111001110001110;
    else if (pixel_index == 5795) oled_data = 16'b1000010001010001;
    else if (pixel_index == 5796 || pixel_index == 5882) oled_data = 16'b1000110001010010;
    else if (pixel_index == 5797) oled_data = 16'b1001110010110011;
    else if (pixel_index == 5800 || pixel_index == 6095) oled_data = 16'b1011010110110110;
    else if (pixel_index == 5803) oled_data = 16'b1010110110111000;
    else if (pixel_index == 5804 || pixel_index == 5900) oled_data = 16'b1010010101110111;
    else if (pixel_index == 5805) oled_data = 16'b1010010011110101;
    else if (pixel_index == 5810) oled_data = 16'b1101011100111010;
    else if (pixel_index == 5815 || pixel_index == 6014) oled_data = 16'b1010110101110101;
    else if (pixel_index == 5856) oled_data = 16'b1000010010110010;
    else if (pixel_index == 5859) oled_data = 16'b1010110101110100;
    else if (pixel_index == 5862 || pixel_index == 5909) oled_data = 16'b1011110111110111;
    else if (pixel_index == 5866) oled_data = 16'b1101011000111001;
    else if (pixel_index == 5867) oled_data = 16'b1101011000111000;
    else if (pixel_index == 5868 || pixel_index == 5997 || pixel_index == 6090) oled_data = 16'b1100111000111000;
    else if (pixel_index == 5870 || pixel_index == 6111) oled_data = 16'b1101111010111001;
    else if (pixel_index == 5878 || pixel_index == 6123) oled_data = 16'b1101011010111001;
    else if (pixel_index == 5879) oled_data = 16'b1100011000110110;
    else if (pixel_index == 5883) oled_data = 16'b0111010000010000;
    else if (pixel_index == 5884) oled_data = 16'b0110001100001100;
    else if ((pixel_index >= 5886) && (pixel_index <= 5887)) oled_data = 16'b0101001010001011;
    else if (pixel_index == 5890) oled_data = 16'b0100101010001011;
    else if (pixel_index == 5891 || pixel_index == 5955 || pixel_index == 5978) oled_data = 16'b0101001010001101;
    else if (pixel_index == 5894) oled_data = 16'b0110101110010000;
    else if ((pixel_index >= 5896) && (pixel_index <= 5897)) oled_data = 16'b1001010010110011;
    else if (pixel_index == 5902 || pixel_index == 6088) oled_data = 16'b1011110111110110;
    else if (pixel_index == 5910) oled_data = 16'b0110001110010001;
    else if (pixel_index == 5911) oled_data = 16'b0100001011001110;
    else if (pixel_index == 5912 || pixel_index == 5992) oled_data = 16'b1000010000010010;
    else if (pixel_index == 5914 || pixel_index == 6124) oled_data = 16'b1100111001111000;
    else if (pixel_index == 5916) oled_data = 16'b1101011001111011;
    else if (pixel_index == 5918) oled_data = 16'b1101011010111000;
    else if (pixel_index == 5954) oled_data = 16'b0111101111001111;
    else if (pixel_index == 5957 || pixel_index == 5974) oled_data = 16'b0111110001010001;
    else if (pixel_index == 5958) oled_data = 16'b0111001111010001;
    else if (pixel_index == 5959) oled_data = 16'b0111001110010001;
    else if (pixel_index == 5961) oled_data = 16'b1000110001010001;
    else if (pixel_index == 5964) oled_data = 16'b1000001110001111;
    else if (pixel_index == 5965) oled_data = 16'b1000001111010000;
    else if (pixel_index == 5966) oled_data = 16'b1000010000010000;
    else if (pixel_index == 5972) oled_data = 16'b1001010001010010;
    else if (pixel_index == 5976 || pixel_index == 6005) oled_data = 16'b0110101101010000;
    else if (pixel_index == 5986 || pixel_index == 6064) oled_data = 16'b0011101000001001;
    else if (pixel_index == 5989) oled_data = 16'b0100101010001101;
    else if (pixel_index == 5993) oled_data = 16'b1001110011110010;
    else if (pixel_index == 5994) oled_data = 16'b1011111000110110;
    else if (pixel_index == 5995) oled_data = 16'b1100111010111001;
    else if (pixel_index == 6002) oled_data = 16'b1011010101110111;
    else if (pixel_index == 6004) oled_data = 16'b1000110010110010;
    else if (pixel_index == 6007) oled_data = 16'b0011101001001101;
    else if (pixel_index == 6009) oled_data = 16'b1011110110110101;
    else if (pixel_index == 6010) oled_data = 16'b1011010111110101;
    else if (pixel_index == 6012) oled_data = 16'b1001010001010100;
    else if (pixel_index == 6013) oled_data = 16'b1010110011110101;
    else if (pixel_index == 6015) oled_data = 16'b1100010111110111;
    else if (pixel_index == 6033) oled_data = 16'b1111111100111110;
    else if (pixel_index == 6035) oled_data = 16'b1110111111111111;
    else if (pixel_index == 6036) oled_data = 16'b1110011111111110;
    else if (pixel_index == 6052 || pixel_index == 6107) oled_data = 16'b0110101101001101;
    else if (pixel_index == 6056) oled_data = 16'b0101101010001100;
    else if (pixel_index == 6058) oled_data = 16'b0111001101001101;
    else if (pixel_index == 6060) oled_data = 16'b0101101100001101;
    else if (pixel_index == 6061) oled_data = 16'b0100101011001101;
    else if (pixel_index == 6065) oled_data = 16'b0011100111001001;
    else if (((pixel_index >= 6066) && (pixel_index <= 6067)) || pixel_index == 6078 || pixel_index == 6080) oled_data = 16'b0010100111001010;
    else if (pixel_index == 6069) oled_data = 16'b0010000110001011;
    else if (pixel_index == 6070) oled_data = 16'b0010100110001010;
    else if (pixel_index == 6071) oled_data = 16'b0011000111001010;
    else if (pixel_index == 6072) oled_data = 16'b0011101000001010;
    else if (pixel_index == 6073) oled_data = 16'b0100001001001010;
    else if (pixel_index == 6074) oled_data = 16'b0010100111001001;
    else if (pixel_index == 6076) oled_data = 16'b0010001000001010;
    else if (pixel_index == 6079) oled_data = 16'b0010000111001001;
    else if (pixel_index == 6081) oled_data = 16'b0011101001001100;
    else if (pixel_index == 6083) oled_data = 16'b0011100110001000;
    else if (pixel_index == 6085) oled_data = 16'b0011001001001101;
    else if (pixel_index == 6086) oled_data = 16'b0100001010001111;
    else if (pixel_index == 6092) oled_data = 16'b1110111100111001;
    else if (pixel_index == 6093) oled_data = 16'b1111011011111011;
    else if (pixel_index == 6097) oled_data = 16'b0110001110010011;
    else if (pixel_index == 6098) oled_data = 16'b1000110000001111;
    else if (pixel_index == 6102) oled_data = 16'b0111001101001111;
    else if (pixel_index == 6104) oled_data = 16'b1001010100110100;
    else if (pixel_index == 6106) oled_data = 16'b0101101011010000;
    else if (pixel_index == 6109) oled_data = 16'b1011010111110110;
    else if (pixel_index == 6113) oled_data = 16'b1110111011111010;
    else if (pixel_index == 6125) oled_data = 16'b1011011000111001;
    else if (pixel_index == 6143) oled_data = 16'b1101111101111111;
    else oled_data = 0;

    end
endmodule
